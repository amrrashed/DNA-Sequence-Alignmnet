
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity ROM_1 is
GENERIC ( bits: INTEGER := 48; -- # of bits per word
 words: INTEGER := 65536); -- # of words in the memory
 PORT ( addr: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 clk:IN STD_LOGIC;
 data: OUT STD_LOGIC_VECTOR (bits-1 DOWNTO 0));
 END ROM_1;

architecture Behavioral of ROM_1 is
TYPE vector_array IS ARRAY (0 TO words-1) OF
 STD_LOGIC_VECTOR (bits-1 DOWNTO 0);
 CONSTANT memory: vector_array := ( 
x"AAAA1111AAAA", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAAA1141AABA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAA1121AACA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAA1121AADA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAA1411ABAA", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"AAAA1441ABBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1421ABCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1421ABDA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1211ACAA", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"AAAA1241ACBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1221ACCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1221ACDA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1211ADAA", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"AAAA1241ADBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1221ADCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAA1221ADDA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"AAAB1111AAAB", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AAAB1121AACB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAB1121AADB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AAAB1411ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AAAB1211ACAB", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"AAAB1221ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAB1221ACDB", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AAAB1211ADAB", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"AAAB1221ADCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAB1221ADDB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA111AAA000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAA111AAA000", 
x"AAAB2111CAAB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAA121ACA000", 
x"AAAB2121CACB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"AAAB2121CADB", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AAAB2211CCAB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"A1A000000000", 
x"AAAB2221CCCB", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAAB2221CCDB", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAAB2211CDAB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"A1A000000000", 
x"AAAB2221CDCB", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAAB2221CDDB", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"AAAB2111DAAB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAA121ACA000", 
x"AAAB2121DACB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"AAAB2121DADB", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AAAB2211DCAB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"A1A000000000", 
x"AAAB2221DCCB", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAAB2221DCDB", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAAB2211DDAB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"A1A000000000", 
x"AAAB2221DDCB", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAAB2221DDDB", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAAC1111AAAC", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAC1141AABC", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAC1121AADC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"AAAC1411ABAC", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAC1441ABBC", 
x"A1A000000000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAC1421ABDC", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AAAC1211ACAC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"AAA121ADA000", 
x"AAAC1211ADAC", 
x"AAA121ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAC1241ADBC", 
x"A1A000000000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAC1221ADDC", 
x"A1A000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AAAC2111CAAC", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"C1C000000000", 
x"AAAC2141CABC", 
x"C1C000000000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAA121ADA000", 
x"C1C000000000", 
x"AAAC2121CADC", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAAC2211CCAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAAC2211CDAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AAAC2111DAAC", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"AAAC2141DABC", 
x"A1A000000000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"AAAC2121DADC", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"AA11AA000000", 
x"AC21DC000000", 
x"AAAC2211DCAC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAAC2211DDAC", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"000000000000", 
x"AAAC2221DDDC", 
x"000000000000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAAD1111AAAD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAD1141AABD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAD1121AACD", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"AAAD1411ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD1441ABBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD1421ABCD", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AA11AA000000", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"AAAD1211ACAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD1241ACBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD1221ACCD", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AA11AA000000", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"AAAD1211ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAA121ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAD2111CAAD", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2141CABD", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2121CACD", 
x"AAA121ADA000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2211CCAD", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAAD2221CCCD", 
x"A1A000000000", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2211CDAD", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAAD2111DAAD", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2141DABD", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2121DACD", 
x"AAA121ADA000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2211DCAD", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAAD2211DDAD", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AABA1141AAAA", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AABA1111AABA", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AABA1141AACA", 
x"AAB121ACB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AABA1141AADA", 
x"AAB121ADB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"AABA1411ABBA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"ABA141ACA000", 
x"ABA141ACA000", 
x"AABA1211ACBA", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AABA1241ACCA", 
x"AAB221CCB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA1241ACDA", 
x"AAB221CDB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"ABA141ADA000", 
x"ABA141ADA000", 
x"AABA1211ADBA", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AABA1241ADCA", 
x"AAB221DCB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA1241ADDA", 
x"AAB221DDB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AAB111AAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"AAB121ACB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AAB121ADB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA211CBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA211DBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AABA2111CABA", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AABA2141CACA", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2141CADA", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"AB11AB000000", 
x"ABA211CBA000", 
x"ABA211CBA000", 
x"BA11BA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2211CCBA", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2211CDBA", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AABA2111DABA", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AABA2141DACA", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2141DADA", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB11AB000000", 
x"ABA211DBA000", 
x"ABA211DBA000", 
x"BA11BA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2211DCBA", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABA2211DDBA", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AABB1111AABB", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AABB1141AACB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AABB1141AADB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AB3B1141ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB3B1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB3B1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"AABB1211ACBB", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"AABB1241ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABB1241ACDB", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"AABB1211ADBB", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"AABB1241ADCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AABB1241ADDB", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"AAB211CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"ABB211CBB000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"ABB211DBB000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AABB2111CABB", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB3B2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB3B2141CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"AABB2211CCBB", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"AABB2211CDBB", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AABB2111DABB", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB3B2141DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB3B2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"AABB2211DCBB", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AABB2211DDBB", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AABC1141AAAC", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AABC1111AABC", 
x"AAB111AAB000", 
x"ABC141AAC000", 
x"AAB121ACB000", 
x"AABC1141AACC", 
x"ABC141AAC000", 
x"AA11AA000000", 
x"AAB121ADB000", 
x"AABC1141AADC", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AABC1411ABBC", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AABC1241ACAC", 
x"C1C000000000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AABC1211ACBC", 
x"AAB121ACB000", 
x"ABC141ACC000", 
x"AAB221CCB000", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"AAB221CDB000", 
x"AABC1241ACDC", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AABC1241ADAC", 
x"A1A000000000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AABC1211ADBC", 
x"AAB121ADB000", 
x"ABC141ADC000", 
x"AAB221DCB000", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AABC1241ADDC", 
x"A1A000000000", 
x"B1B000000000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"B1B000000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AABC2141CAAC", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AABC2111CABC", 
x"AAB211CAB000", 
x"C1C000000000", 
x"AAB121ACB000", 
x"AABC2141CACC", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB121ADB000", 
x"AABC2141CADC", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AABC2211CCBC", 
x"AAB221CCB000", 
x"C1C000000000", 
x"AAB221CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AABC2211CDBC", 
x"AAB221CDB000", 
x"C1C000000000", 
x"AAB221DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221DDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AABC2141DAAC", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AABC2111DABC", 
x"AAB211DAB000", 
x"C1C000000000", 
x"AAB121ACB000", 
x"AABC2141DACC", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"AABC2141DADC", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AABC2211DCBC", 
x"AAB221DCB000", 
x"C1C000000000", 
x"AAB221CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAB221CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AABC2211DDBC", 
x"AAB221DDB000", 
x"C1C000000000", 
x"AAB221DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"C1C000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AABD1141AAAD", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AABD1111AABD", 
x"AA11AA000000", 
x"AAB121ACB000", 
x"AA11AA000000", 
x"AABD1141AACD", 
x"AA11AA000000", 
x"AAB121ADB000", 
x"AA11AA000000", 
x"AABD1141AADD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AABD1411ABBD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"AABD1241ACAD", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AABD1211ACBD", 
x"A1A000000000", 
x"AAB221CCB000", 
x"A1A000000000", 
x"AABD1241ACCD", 
x"ABD141ACD000", 
x"AAB221CDB000", 
x"ABD141ACD000", 
x"AABD1241ACDD", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"AABD1241ADAD", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AABD1211ADBD", 
x"A1A000000000", 
x"AAB221DCB000", 
x"A1A000000000", 
x"AABD1241ADCD", 
x"ABD141ADD000", 
x"AAB221DDB000", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"B1B000000000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"B1B000000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"AAB211CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AAB211DAB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AABD2111CABD", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"AABD2141CACD", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"AABD2141CADD", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AABD2211CCBD", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AABD2211CDBD", 
x"A1A000000000", 
x"AAB221DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AABD2111DABD", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"AABD2141DACD", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"AABD2141DADD", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AABD2211DCBD", 
x"A1A000000000", 
x"AAB221CCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AAB221CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AABD2211DDBD", 
x"A1A000000000", 
x"AAB221DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AACA1121AAAA", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AACA1141AABA", 
x"AA11AA000000", 
x"AAC141ABC000", 
x"AA11AA000000", 
x"AACA1111AACA", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AACA1141AADA", 
x"AA11AA000000", 
x"AAC121ADC000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ACA141ABA000", 
x"AC11AC000000", 
x"ACA141ABA000", 
x"AACA1441ABBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AACA1411ABCA", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AACA1441ABDA", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AACA1211ACCA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"ACA141ADA000", 
x"AAC211DAC000", 
x"ACA141ADA000", 
x"AACA1241ADBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AACA1211ADCA", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AACA1241ADDA", 
x"A1A000000000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAC211CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAC111AAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AACA2111CACA", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAC121ADC000", 
x"CA11CA000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"ACA211CCA000", 
x"AAC211CAC000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AACA2211CCCA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211DAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AACA2211CDCA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AACA2141DABA", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"AACA2111DACA", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AACA2141DADA", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACA211DCA000", 
x"ACA211DCA000", 
x"AAC211CAC000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AACA2211DCCA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AACA2211DDCA", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AA11AA000000", 
x"AACB1121AAAB", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"ACB121AAB000", 
x"AACB1141AABB", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"AAC111AAC000", 
x"AACB1111AACB", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AACB1141AADB", 
x"AAC121ADC000", 
x"AA11AA000000", 
x"CB21AB000000", 
x"AACB1421ABAB", 
x"AC11AC000000", 
x"CB21AB000000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"CB21AB000000", 
x"AACB1411ABCB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AACB1441ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"AACB1221ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AACB1211ACCB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"AACB1221ADAB", 
x"AAC211DAC000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"AAC121ADC000", 
x"AACB1211ADCB", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AACB1241ADDB", 
x"AAC221DDC000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACB121AAB000", 
x"AAC111AAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"AAC121ADC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC211CAC000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"ACB211CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB211DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AACB2121CAAB", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"ACB221CAB000", 
x"AACB2141CABB", 
x"ACB221CAB000", 
x"ACB221CAB000", 
x"AAC211CAC000", 
x"AACB2111CACB", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"AACB2141CADB", 
x"AAC121ADC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"AA11AA000000", 
x"AACB2221CCAB", 
x"AAC211CAC000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"AACB2211CCCB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AACB2221CDAB", 
x"AAC211DAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AACB2211CDCB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AACB2121DAAB", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"ACB221DAB000", 
x"AACB2141DABB", 
x"ACB221DAB000", 
x"ACB221DAB000", 
x"AAC211DAC000", 
x"AACB2111DACB", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"AACB2141DADB", 
x"AAC121ADC000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AACB2221DCAB", 
x"AAC211CAC000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AACB2211DCCB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"AACB2221DDAB", 
x"AAC211DAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"AACB2211DDCB", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AACC1141AABC", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AACC1111AACC", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AACC1141AADC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AACC1441ABBC", 
x"A1A000000000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AACC1411ABCC", 
x"AAC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AACC1441ABDC", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AACC1241ADBC", 
x"A1A000000000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AACC1211ADCC", 
x"AAC121ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AACC1241ADDC", 
x"A1A000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAC141ABC000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AACC2111CACC", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAC121ADC000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211DAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AACC2211CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AACC2111DACC", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"AA11AA000000", 
x"AC21DC000000", 
x"AAC211CAC000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AACC2211DDCC", 
x"AAC221DDC000", 
x"A1A000000000", 
x"000000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AACD1121AAAD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC141ABC000", 
x"AACD1141AABD", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AACD1111AACD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC121ADC000", 
x"AACD1141AADD", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AACD1421ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AACD1441ABBD", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AACD1411ABCD", 
x"ACD141ABD000", 
x"ACD141ABD000", 
x"AC21DC000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AACD1211ACCD", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"AACD1221ADAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AACD1241ADBD", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AACD1211ADCD", 
x"ACD141ADD000", 
x"ACD141ADD000", 
x"AAC221DDC000", 
x"ACD141ADD000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"ACD141ADD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"AAC221DDC000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAC141ABC000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AACD2111CACD", 
x"C1C000000000", 
x"C1C000000000", 
x"AAC121ADC000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AACD2211CCCD", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AAC211DAC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"AACD2141DABD", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AACD2111DACD", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"AACD2141DADD", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AC21DC000000", 
x"AAC211CAC000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AACD2211DCCD", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"AACD2211DDCD", 
x"A1A000000000", 
x"D1D000000000", 
x"AAC221DDC000", 
x"D1D000000000", 
x"AADA1121AAAA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AADA1141AABA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADA1141AACA", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADA1111AADA", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"AD11AD000000", 
x"AADA1441ABBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADA1441ABCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADA1411ABDA", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AA11AA000000", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"AAD211CAD000", 
x"AADA1241ACBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADA1241ACCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADA1211ACDA", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AADA1211ADDA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"ADA211CDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AA11AA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AADA2141CABA", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"AADA2141CACA", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AADA2111CADA", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"AADA2211CCDA", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AA11AA000000", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AADA2211CDDA", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AAD121ACD000", 
x"AADA2111DADA", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AADA2211DCDA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AADA2211DDDA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AADB1121AAAB", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"ADB121AAB000", 
x"AADB1141AABB", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"AA11AA000000", 
x"AADB1141AACB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AADB1111AADB", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"DB21AB000000", 
x"AADB1421ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"DB21AB000000", 
x"AADB1441ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AADB1411ABDB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AA11AA000000", 
x"AADB1221ACAB", 
x"A1A000000000", 
x"AAD211CAD000", 
x"ADB141ACB000", 
x"AADB1241ACBB", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"AADB1241ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AADB1211ACDB", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AA11AA000000", 
x"AADB1221ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AADB1241ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AADB1211ADDB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"AAD111AAD000", 
x"B1B000000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AADB2121CAAB", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"ADB221CAB000", 
x"AADB2141CABB", 
x"ADB221CAB000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AADB2141CACB", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211CAD000", 
x"AADB2111CADB", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AADB2221CCAB", 
x"A1A000000000", 
x"AAD211CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"A1A000000000", 
x"AADB2211CCDB", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AA11AA000000", 
x"AADB2221CDAB", 
x"A1A000000000", 
x"AAD211DAD000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AADB2211CDDB", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AA11AA000000", 
x"AADB2121DAAB", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"ADB221DAB000", 
x"AADB2141DABB", 
x"ADB221DAB000", 
x"ADB221DAB000", 
x"A1A000000000", 
x"AADB2141DACB", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211DAD000", 
x"AADB2111DADB", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AA11AA000000", 
x"AADB2221DCAB", 
x"A1A000000000", 
x"AAD211CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AADB2211DCDB", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AADB2221DDAB", 
x"A1A000000000", 
x"AAD211DAD000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AADB2211DDDB", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADC1121AAAC", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADC1141AABC", 
x"AA11AA000000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"AADC1141AACC", 
x"ADC121AAC000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AADC1111AADC", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AADC1421ABAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADC1441ABBC", 
x"A1A000000000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AADC1411ABDC", 
x"AAD141ABD000", 
x"AA11AA000000", 
x"DC21AC000000", 
x"AADC1221ACAC", 
x"AAD211CAD000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"AADC1241ACBC", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AADC1211ACDC", 
x"AAD121ACD000", 
x"AA11AA000000", 
x"AD11AD000000", 
x"AADC1221ADAC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AADC1241ADBC", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AADC1211ADDC", 
x"AD11AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ADC121AAC000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"AAD141ABD000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"AAD121ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD211CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"ADC221DAC000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADC2121CAAC", 
x"AAD111AAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AADC2141CABC", 
x"AAD141ABD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AADC2141CACC", 
x"AAD121ACD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AADC2111CADC", 
x"AAD211CAD000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD211CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AADC2211CCDC", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD211DAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"AADC2211CDDC", 
x"C1C000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADC2121DAAC", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADC2141DABC", 
x"AAD141ABD000", 
x"ADC221DAC000", 
x"ADC221DAC000", 
x"AADC2141DACC", 
x"AAD121ACD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AADC2111DADC", 
x"AAD211DAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AADC2221DDAC", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"A1A000000000", 
x"D1D000000000", 
x"AADC2211DDDC", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADD1141AABD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AADD1141AACD", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AADD1111AADD", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADD1441ABBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADD1441ABCD", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AADD1411ABDD", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADD1241ACBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AADD1241ACCD", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AADD1211ACDD", 
x"AA11AA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AADD2111CADD", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"A1A000000000", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AADD2211CCDD", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AADD2111DADD", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AADD2211DCDD", 
x"AA11AA000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AAD211DAD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ABAA1411AAAA", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ABAA1111ABAA", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABAA1141ABBA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAA1121ABCA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAA1121ABDA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAA1411ACAA", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABA141ACA000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAA1421ACCA", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAA1421ACDA", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAA1411ADAA", 
x"AB11AB000000", 
x"ABA141ADA000", 
x"ABA141ADA000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAA1421ADCA", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAA1421ADDA", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"AB11AB000000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"ABA211CBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"AB11AB000000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"ABA211DBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAA2111CBAA", 
x"AB11AB000000", 
x"ABA211CBA000", 
x"ABA211CBA000", 
x"BA11BA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAA2121CBCA", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAA2121CBDA", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAA2111DBAA", 
x"AB11AB000000", 
x"ABA211DBA000", 
x"ABA211DBA000", 
x"BA11BA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAA2121DBCA", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAA2121DBDA", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"ABA141AAA000", 
x"ABAB1411AAAB", 
x"ABA141AAA000", 
x"ABA141AAA000", 
x"ABA111ABA000", 
x"ABAB1141AB3B", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABAB1421AACB", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"ABAB1421AADB", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"ABAB1111ABAB", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABAB1141AB3B", 
x"ABAB1141ABBB", 
x"ABAB1141AB3B", 
x"ABAB1141AB3B", 
x"AB11AB000000", 
x"ABAB1121ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAB1121ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABAB1411ACAB", 
x"ABA141ACA000", 
x"ABA141ACA000", 
x"ABA211CBA000", 
x"ABAB2141CB3B", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABAB1421ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAB1421ACDB", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"ABAB1411ADAB", 
x"ABA141ADA000", 
x"ABA141ADA000", 
x"ABA211DBA000", 
x"ABAB2141DB3B", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ABAB1421ADCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABAB1421ADDB", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3AB1411BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA3B1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA3B1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB121BCB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB121BDB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B3AB1411BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B3AB1421BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1421BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1411BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B3AB1421BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1421BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"ABAB1141AB3B", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"ABAB2111CBAB", 
x"ABA211CBA000", 
x"ABA211CBA000", 
x"BA11BA000000", 
x"ABAB2141CBBB", 
x"ABAB2141CB3B", 
x"ABAB2141CB3B", 
x"AB21CB000000", 
x"ABAB2121CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAB2121CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"ABAB2141CB3B", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"ABAB2141DB3B", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"ABAB1141AB3B", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"ABAB2111DBAB", 
x"ABA211DBA000", 
x"ABA211DBA000", 
x"BA11BA000000", 
x"ABAB2141DBBB", 
x"ABAB2141DB3B", 
x"ABAB2141DB3B", 
x"AB21DB000000", 
x"ABAB2121DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAB2121DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211CBA000", 
x"ABAB2141CB3B", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"ABAB2141DB3B", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"ABAC1411AAAC", 
x"ABA141AAA000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB21CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"ABAC1421AADC", 
x"A1A000000000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABAC1111ABAC", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAC1141ABBC", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAC1121ABCC", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAC1121ABDC", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB11AB000000", 
x"ABAC1411ACAC", 
x"AC11AC000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AC11AC000000", 
x"AB21CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AB21DB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ABA141ADA000", 
x"AB11AB000000", 
x"ABAC1411ADAC", 
x"ABA141ADA000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"AB21CB000000", 
x"ABAC1421ADCC", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABAC1421ADDC", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"BAC141BBC000", 
x"BAC121BCC000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B3AC1411BCAC", 
x"B1B000000000", 
x"ABA211CBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B3AC1411BDAC", 
x"B1B000000000", 
x"ABA211DBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB21CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABA211CBA000", 
x"AB11AB000000", 
x"ABAC2111CBAC", 
x"ABA211CBA000", 
x"BA11BA000000", 
x"AB21CB000000", 
x"ABAC2141CBBC", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAC2121CBCC", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAC2121CBDC", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB21CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ABA141ADA000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB11AB000000", 
x"ABAC2111DBAC", 
x"ABA211DBA000", 
x"BA11BA000000", 
x"AB21DB000000", 
x"ABAC2141DBBC", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAC2121DBCC", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAC2121DBDC", 
x"AB21DB000000", 
x"AC21DC000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AC21DC000000", 
x"AB21CB000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"AB21CB000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"000000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"ABA141AAA000", 
x"ABAD1411AAAD", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABAD1421AACD", 
x"AD11AD000000", 
x"AB21DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABAD1111ABAD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAD1141ABBD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAD1121ABCD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABAD1121ABDD", 
x"ABA141ACA000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABAD1411ACAD", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABAD1421ACCD", 
x"A1A000000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ABAD1421ACDD", 
x"AD11AD000000", 
x"AB11AB000000", 
x"AD11AD000000", 
x"ABAD1411ADAD", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AD11AD000000", 
x"AB21CB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AB21DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD121BDD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B3AD1411BCAD", 
x"ABA211CBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B3AD1411BDAD", 
x"ABA211DBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"AB21DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ABA211CBA000", 
x"AB11AB000000", 
x"ABA211CBA000", 
x"ABAD2111CBAD", 
x"BA11BA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAD2141CBBD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAD2121CBCD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABAD2121CBDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"AB21DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ABA211DBA000", 
x"AB11AB000000", 
x"ABA211DBA000", 
x"ABAD2111DBAD", 
x"BA11BA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAD2141DBBD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAD2121DBCD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABAD2121DBDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ABBA1441AAAA", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1411AABA", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABBA1441AACA", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1441AADA", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1141ABAA", 
x"AB3B1141ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABBA1111ABBA", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABBA1141ABCA", 
x"AB3B1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABBA1141ABDA", 
x"AB3B1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABBA1441ACAA", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1411ACBA", 
x"ABB211CBB000", 
x"ABB141ACB000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1441ACDA", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1441ADAA", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1411ADBA", 
x"ABB211DBB000", 
x"ABB141ADB000", 
x"ABB141ADB000", 
x"ABBA1441ADCA", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBA1441ADDA", 
x"AB21DB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B3BA1411BABA", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"AB11AB000000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"B3BA1411BCBA", 
x"ABB211CBB000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"AB11AB000000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"B3BA1411BDBA", 
x"ABB211DBB000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABBA2111CBBA", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABBA2141CBCA", 
x"AB3B2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABBA2141CBDA", 
x"AB3B2141CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABBA2111DBBA", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABBA2141DBCA", 
x"AB3B2141DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABBA2141DBDA", 
x"AB3B2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABBB1141ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABBB1111ABBB", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"ABBB1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABBB1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"ABBB1411ACBB", 
x"ABB141ACB000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBB1441ACDB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"ABBB1411ADBB", 
x"ABB141ADB000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"ABBB1441ADCB", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABBB1441ADDB", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"ABB111ABB000", 
x"BBB141BAB000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BB3B1441BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB3B1141BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB3B1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB3B1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B3BB1411BCBB", 
x"BBB141BCB000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B3BB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3BB1441BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B3BB1411BDBB", 
x"BBB141BDB000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"BB3B1441BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3BB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABBB2141CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"ABBB2111CBBB", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"ABBB2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABBB2141CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABBB2141DBAB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"ABBB2111DBBB", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"ABBB2141DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABBB2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABBC1441AAAC", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABBC1411AABC", 
x"AB11AB000000", 
x"C1C000000000", 
x"ABB141ACB000", 
x"ABBC1441AACC", 
x"C1C000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"ABBC1441AADC", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB3B1141ABAB", 
x"ABBC1141ABAC", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABBC1111ABBC", 
x"ABB111ABB000", 
x"BC11BC000000", 
x"AB3B1141ABCB", 
x"ABBC1141ABCC", 
x"BC11BC000000", 
x"AB11AB000000", 
x"AB3B1141ABDB", 
x"ABBC1141ABDC", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABBC1441ACAC", 
x"C1C000000000", 
x"ABB141ACB000", 
x"ABB211CBB000", 
x"ABBC1411ACBC", 
x"ABB141ACB000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABBC1441ACDC", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABBC1441ADAC", 
x"A1A000000000", 
x"ABB141ADB000", 
x"ABB211DBB000", 
x"ABBC1411ADBC", 
x"ABB141ADB000", 
x"C1C000000000", 
x"AB21CB000000", 
x"ABBC1441ADCC", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABBC1441ADDC", 
x"A1A000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"B3BC1411BABC", 
x"AB11AB000000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"ABB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"ABB211CBB000", 
x"B3BC1411BCBC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"ABB211DBB000", 
x"B3BC1411BDBC", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"ABB141ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"ABBC2141CBAC", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABBC2111CBBC", 
x"ABB211CBB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"AB3B2141CBDB", 
x"ABBC2141CBDC", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"ABB141ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"ABBC2141DBAC", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABBC2111DBBC", 
x"ABB211DBB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"AB3B2141DBDB", 
x"ABBC2141DBDC", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABBD1441AAAD", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"ABBD1411AABD", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"ABBD1441AACD", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"ABBD1441AADD", 
x"AB11AB000000", 
x"AB3B1141ABAB", 
x"AB11AB000000", 
x"ABBD1141ABAD", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABBD1111ABBD", 
x"AB11AB000000", 
x"AB3B1141ABCB", 
x"AB11AB000000", 
x"ABBD1141ABCD", 
x"AB11AB000000", 
x"AB3B1141ABDB", 
x"AB11AB000000", 
x"ABBD1141ABDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABBD1441ACAD", 
x"ABB141ACB000", 
x"ABB211CBB000", 
x"ABB141ACB000", 
x"ABBD1411ACBD", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ABBD1441ACDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABBD1441ADAD", 
x"ABB141ADB000", 
x"ABB211DBB000", 
x"ABB141ADB000", 
x"ABBD1411ADBD", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABBD1441ADCD", 
x"A1A000000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ABBD1441ADDD", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"B3BD1411BABD", 
x"B1B000000000", 
x"ABB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"ABB141ADB000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"ABB211CBB000", 
x"B3B141BCB000", 
x"B3BD1411BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"ABB211DBB000", 
x"B3B141BDB000", 
x"B3BD1411BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"ABBD2141CBAD", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABBD2111CBBD", 
x"AB21CB000000", 
x"AB3B2141CBCB", 
x"AB21CB000000", 
x"ABBD2141CBCD", 
x"BD11BD000000", 
x"AB3B2141CBDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"ABBD2141DBAD", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABBD2111DBBD", 
x"AB21DB000000", 
x"AB3B2141DBCB", 
x"AB21DB000000", 
x"ABBD2141DBCD", 
x"BD11BD000000", 
x"AB3B2141DBDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ABCA1421AAAA", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABCA1411AACA", 
x"AB21CB000000", 
x"ABC141AAC000", 
x"ABC141AAC000", 
x"ABCA1441AADA", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"ABCA1121ABAA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCA1141ABBA", 
x"AB11AB000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"ABCA1111ABCA", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABCA1141ABDA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"ABCA1411ACCA", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABCA1421ADAA", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"ABCA1411ADCA", 
x"AB21CB000000", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"ABCA1441ADDA", 
x"AB21DB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"AB11AB000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"B3CA1411BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA121BAA000", 
x"AB11AB000000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"AB11AB000000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"B3CA1411BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ABCA2121CBAA", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABCA2141CBBA", 
x"AB21CB000000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"ABCA2111CBCA", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABCA2141CBDA", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"ABCA2121DBAA", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABCA2141DBBA", 
x"AB21DB000000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"ABCA2111DBCA", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABCA2141DBDA", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABCB1141AB3B", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"ABCB1411AACB", 
x"ABC141AAC000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"ABCB1441AADB", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABCB1121ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCB1141AB3B", 
x"ABCB1141ABBB", 
x"ABCB1141AB3B", 
x"ABCB1141AB3B", 
x"ABC111ABC000", 
x"ABCB1111ABCB", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABCB1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ABC211CBC000", 
x"CB11CB000000", 
x"ABC141ACC000", 
x"ABCB1411ACCB", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABCB2141DB3B", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"ABCB1411ADCB", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"ABCB1441ADDB", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"ABC111ABC000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC3B1241BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB121BAB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BCB141BDB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"B3CB1411BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABCB1141AB3B", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"ABCB2121CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ABCB2141CBBB", 
x"BC11BC000000", 
x"CB11CB000000", 
x"ABC211CBC000", 
x"ABCB2111CBCB", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"CB11CB000000", 
x"ABCB2141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ABC211CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABCB2141DB3B", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABCB1141AB3B", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABCB2121DBAB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABCB2141DB3B", 
x"ABCB2141DBBB", 
x"BC11BC000000", 
x"ABCB2141DB3B", 
x"ABC211DBC000", 
x"ABCB2111DBCB", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"ABCB2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ABC211CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABCB2141DB3B", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"AB21CB000000", 
x"ABCC1411AACC", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCC1121ABAC", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCC1141ABBC", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABCC1111ABCC", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCC1141ABDC", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABCC1421ACAC", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"ABCC1411ACCC", 
x"CC11CC000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABCC1421ADAC", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"AB21CB000000", 
x"ABCC1411ADCC", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABCC1441ADDC", 
x"A1A000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"BCC141BDC000", 
x"B3CC1411BDCC", 
x"BCC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"ABCC2121CBAC", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABCC2111CBCC", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABCC2141CBDC", 
x"AB21CB000000", 
x"CC11CC000000", 
x"AB11AB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"ABC211CBC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"ABCC2121DBAC", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABCC2111DBCC", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABCC2141DBDC", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"ABCD1421AAAD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"AB21CB000000", 
x"ABC141AAC000", 
x"ABCD1411AACD", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"ABCD1441AADD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCD1121ABAD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BC11BC000000", 
x"ABCD1141ABBD", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABCD1111ABCD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABCD1141ABDD", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"ABCD1411ACCD", 
x"CD11CD000000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"ABCD1421ADAD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"AB21CB000000", 
x"ABC141ADC000", 
x"ABCD1411ADCD", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"ABCD1441ADDD", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BDD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"CD11CD000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"ABCD2121CBAD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BC11BC000000", 
x"ABCD2141CBBD", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABCD2111CBCD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABCD2141CBDD", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AB11AB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"AB21CB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"ABCD2121DBAD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BC11BC000000", 
x"ABCD2141DBBD", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABCD2111DBCD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABCD2141DBDD", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ABDA1421AAAA", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABDA1441AACA", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"ABDA1411AADA", 
x"AB21DB000000", 
x"ABD141AAD000", 
x"ABD141AAD000", 
x"ABDA1121ABAA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDA1141ABBA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDA1141ABCA", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDA1111ABDA", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABDA1421ACAA", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABDA1411ACDA", 
x"AB21DB000000", 
x"ABD141ACD000", 
x"ABD141ACD000", 
x"DA11DA000000", 
x"AB11AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"ABDA1441ADCA", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABDA1411ADDA", 
x"AB21DB000000", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"BDA121BAA000", 
x"AB11AB000000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA121BAA000", 
x"AB11AB000000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"AB11AB000000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"ABDA2121CBAA", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDA2141CBBA", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"ABDA2141CBCA", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDA2111CBDA", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB11AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB11AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"DA11DA000000", 
x"AB21CB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ABDA2121DBAA", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABDA2141DBBA", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"ABDA2141DBCA", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABDA2111DBDA", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB11AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"ABDB1141AB3B", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"ABDB1441AACB", 
x"A1A000000000", 
x"ABD141ACD000", 
x"ABD141AAD000", 
x"ABDB1411AADB", 
x"ABD141AAD000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"ABDB1121ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDB1141AB3B", 
x"ABDB1141ABBB", 
x"ABDB1141AB3B", 
x"ABDB1141AB3B", 
x"AB11AB000000", 
x"ABDB1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABDB1111ABDB", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABDB2141CB3B", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"ABDB1411ACDB", 
x"ABD141ACD000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"ABDB1441ADCB", 
x"A1A000000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"ABDB1411ADDB", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BD3B1241BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB121BAB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDB141BCB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B3DB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD3B1141BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD3B1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3DB1411BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"ABDB1141AB3B", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"DB11DB000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"AB21CB000000", 
x"ABDB2121CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDB2141CB3B", 
x"ABDB2141CBBB", 
x"ABDB2141CB3B", 
x"BD11BD000000", 
x"AB21CB000000", 
x"ABDB2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"ABDB2111CBDB", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABDB2141CB3B", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"ABDB1141AB3B", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"DB11DB000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"DB11DB000000", 
x"ABDB2121DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"ABDB2141DBBB", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"ABDB2141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"ABD211DBD000", 
x"ABDB2111DBDB", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"ABDB2141CB3B", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABDC1421AAAC", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"DC21AC000000", 
x"AB21CB000000", 
x"ABDC1441AACC", 
x"DC21AC000000", 
x"ABD141AAD000", 
x"AB21DB000000", 
x"ABDC1411AADC", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDC1121ABAC", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDC1141ABBC", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDC1141ABCC", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABDC1111ABDC", 
x"ABD111ABD000", 
x"DC21AC000000", 
x"AB11AB000000", 
x"ABDC1421ACAC", 
x"DC21AC000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"DC21AC000000", 
x"AB21CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"AB21DB000000", 
x"ABDC1411ACDC", 
x"DC21AC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABDC1421ADAC", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ABD141ADD000", 
x"AB21DB000000", 
x"ABDC1411ADDC", 
x"ABD141ADD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BD11BD000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"ABD141ADD000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"ABDC2121CBAC", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDC2141CBBC", 
x"BD11BD000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDC2141CBCC", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABDC2111CBDC", 
x"ABD211CBD000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"DC21AC000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"DC21AC000000", 
x"AB21CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"ABD141ADD000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"ABDC2121DBAC", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABDC2141DBBC", 
x"BD11BD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABDC2141DBCC", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABDC2111DBDC", 
x"ABD211DBD000", 
x"DC11DC000000", 
x"AB11AB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"DC21AC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"ABD141AAD000", 
x"AB21DB000000", 
x"ABD141AAD000", 
x"ABDD1411AADD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDD1121ABAD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDD1141ABBD", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABDD1141ABCD", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABDD1111ABDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABDD1421ACAD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"AB21DB000000", 
x"ABD141ACD000", 
x"ABDD1411ACDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABDD1421ADAD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABDD1441ADCD", 
x"DD11DD000000", 
x"AB21DB000000", 
x"DD11DD000000", 
x"ABDD1411ADDD", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"DD11DD000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"ABDD2121CBAD", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABDD2141CBCD", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABDD2111CBDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AB21DB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"DD11DD000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"ABDD2121DBAD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABDD2141DBCD", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABDD2111DBDD", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AB11AB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"DD11DD000000", 
x"AB21CB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AB21DB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ACAA1211AAAA", 
x"ACA121AAA000", 
x"AC11AC000000", 
x"ACA121AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ACAA1411ABAA", 
x"ACA141ABA000", 
x"AC11AC000000", 
x"ACA141ABA000", 
x"ACAA1441ABBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAA1421ABDA", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACAA1111ACAA", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACAA1141ACBA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAA1121ACCA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAA1121ACDA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAA1411ADAA", 
x"ACA141ADA000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACAA1441ADBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAA1421ADDA", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACA121AAA000", 
x"AA11AA000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"AC11AC000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAA2111CCAA", 
x"ACA211CCA000", 
x"AC11AC000000", 
x"ACA211CCA000", 
x"ACAA2141CCBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAA2121CCDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"AC11AC000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211DCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA121AAA000", 
x"AA11AA000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACAA2111DCAA", 
x"ACA211DCA000", 
x"AC11AC000000", 
x"ACA211DCA000", 
x"ACAA2141DCBA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACA211CCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAA2121DCDA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACA121AAA000", 
x"ACAB1211AAAB", 
x"AC11AC000000", 
x"ACA121AAA000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"ACA111ACA000", 
x"ACAB1221AACB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACAB1221AADB", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ACAB1411ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ACA111ACA000", 
x"ACAB1111ACAB", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACAB1141AC3B", 
x"ACAB1141ACBB", 
x"ACAB1141AC3B", 
x"ACAB1141AC3B", 
x"AC11AC000000", 
x"ACAB1121ACCB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAB1121ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACAB1411ADAB", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"CAB221ADB000", 
x"ACAB1441ADBB", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"ACA211DCA000", 
x"ACAB1421ADCB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACAB1421ADDB", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ACA111ACA000", 
x"ACAB1141AC3B", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211CCA000", 
x"CAB121CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211DCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"ACAB2211CAAB", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"ACA111ACA000", 
x"ACAB1141AC3B", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA3B1141CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ACA211CCA000", 
x"ACAB2111CCAB", 
x"AC11AC000000", 
x"ACA211CCA000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"ACA211CCA000", 
x"ACAB2121CCCB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAB2121CCDB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"ACA211DCA000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA121AAA000", 
x"ACAB2211DAAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ACA111ACA000", 
x"ACAB1141AC3B", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACAB2221DADB", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ACA211DCA000", 
x"ACAB2111DCAB", 
x"AC11AC000000", 
x"ACA211DCA000", 
x"AB21CB000000", 
x"ACAB2141DCBB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ACA211CCA000", 
x"ACAB2121DCCB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAB2121DCDB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ACA211DCA000", 
x"AB21CB000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACA121AAA000", 
x"ACA121AAA000", 
x"ACAC1211AAAC", 
x"ACA121AAA000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"ACAC1241AABC", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"ACAC1221AADC", 
x"A1A000000000", 
x"ACA141ABA000", 
x"ACA141ABA000", 
x"ACAC1411ABAC", 
x"ACA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACAC1441ABBC", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ACAC1421ABCC", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACAC1421ABDC", 
x"A1A000000000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACAC1111ACAC", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAC1141ACBC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAC1121ACCC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAC1121ACDC", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACA141ADA000", 
x"ACAC1411ADAC", 
x"ACA141ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACAC1441ADBC", 
x"A1A000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"ACAC1421ADCC", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACAC1421ADDC", 
x"A1A000000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"ACA211CCA000", 
x"ACAC2111CCAC", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAC2141CCBC", 
x"C1C000000000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAC2121CCDC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACA211DCA000", 
x"ACA211DCA000", 
x"ACAC2111DCAC", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAC2141DCBC", 
x"AC21DC000000", 
x"ACA211CCA000", 
x"AC21DC000000", 
x"ACAC2121DCCC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAC2121DCDC", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"ACA121AAA000", 
x"ACA121AAA000", 
x"AC11AC000000", 
x"ACAD1211AAAD", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACAD1241AABD", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"ACA141ABA000", 
x"ACA141ABA000", 
x"AC11AC000000", 
x"ACAD1411ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACAD1441ABBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"ACAD1421ABDD", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACAD1111ACAD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAD1141ACBD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAD1121ACCD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACAD1121ACDD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AC11AC000000", 
x"ACAD1411ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ACA211DCA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"AC11AC000000", 
x"CAD211AAD000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"ACA211CCA000", 
x"ACA211CCA000", 
x"AC11AC000000", 
x"ACAD2111CCAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAD2141CCBD", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACAD2121CCCD", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211DCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACAD2211DAAD", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACA211DCA000", 
x"ACA211DCA000", 
x"AC11AC000000", 
x"ACAD2111DCAD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAD2141DCBD", 
x"ACA211CCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAD2121DCCD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACAD2121DCDD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACBA1241AAAA", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACBA1211AABA", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACBA1241AADA", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"ACBA1411ABBA", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"ACBA1141ACAA", 
x"AC3B1141ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACBA1111ACBA", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACBA1141ACCA", 
x"ACB211CCB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACBA1141ACDA", 
x"AC3B1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACBA1441ADAA", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACBA1411ADBA", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACBA1441ADDA", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ACB121AAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ACB111ACB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"ACB211CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB211DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"CBA141CAA000", 
x"ACBA2211CABA", 
x"ACB141ABB000", 
x"ACB221CAB000", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ACBA2141CCAA", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"CBA141CCA000", 
x"ACBA2111CCBA", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACBA2141CCCA", 
x"ACB211CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACBA2141CCDA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB211DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACBA2211DABA", 
x"ACB141ABB000", 
x"ACB221DAB000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACBA2141DCAA", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ACBA2111DCBA", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACBA2141DCCA", 
x"ACB211CCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACBA2141DCDA", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"ACBB1211AABB", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACBB1241AADB", 
x"AC21DC000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB3B2141ABAB", 
x"AC11AC000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"ACBB1411ABBB", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB3B2141ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"ACBB1141ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"ACBB1111ACBB", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"ACBB1141ACCB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACBB1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACBB1441ADAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"ACBB1411ADBB", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACBB1441ADDB", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"CBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CBB141CAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"ACB211CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"ACB211DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"ACBB2211CABB", 
x"CBB141CAB000", 
x"CBB141CAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB3B1141CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB3B1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"ACBB2141CCAB", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"ACBB2111CCBB", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACBB2141CCDB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"BB11BB000000", 
x"CBB141CDB000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"ACB211DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"ACBB2211DABB", 
x"ACB221DAB000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACBB2141DCAB", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"ACBB2111DCBB", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"ACB211CCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACBB2141DCDB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACBC1211AABC", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"ACBC1241AADC", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB21AB000000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACBC1411ABBC", 
x"ACB141ABB000", 
x"CBC211ABC000", 
x"CB11CB000000", 
x"CBC211ABC000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"AC3B1141ACAB", 
x"ACBC1141ACAC", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACBC1111ACBC", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"ACB211CCB000", 
x"ACBC1141ACCC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"ACBC1141ACDC", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACBC1411ADBC", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACBC1441ADDC", 
x"A1A000000000", 
x"B1B000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB141ABB000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"ACB211CCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB211DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"ACB141ABB000", 
x"ACBC2211CABC", 
x"ACB221CAB000", 
x"CBC141CAC000", 
x"ACB111ACB000", 
x"CBC141CAC000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"ACBC2141CCAC", 
x"C1C000000000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACBC2111CCBC", 
x"ACB211CCB000", 
x"CBC141CCC000", 
x"ACB211CCB000", 
x"CBC141CCC000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"B1B000000000", 
x"ACBC2141CCDC", 
x"C1C000000000", 
x"C1C000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"ACB211DCB000", 
x"CBC141CDC000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"ACB141ABB000", 
x"ACBC2211DABC", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACB221CAB000", 
x"ACBC2141DCAC", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACBC2111DCBC", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"ACB211CCB000", 
x"ACBC2141DCCC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"ACBC2141DCDC", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"ACBD1241AAAD", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACBD1211AABD", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"ACBD1241AADD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB21AB000000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACBD1411ABBD", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"AC11AC000000", 
x"AC3B1141ACAB", 
x"AC11AC000000", 
x"ACBD1141ACAD", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACBD1111ACBD", 
x"AC11AC000000", 
x"ACB211CCB000", 
x"AC11AC000000", 
x"ACBD1141ACCD", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"AC11AC000000", 
x"ACBD1141ACDD", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"ACBD1441ADAD", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACBD1411ADBD", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACBD1441ADDD", 
x"B1B000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"B1B000000000", 
x"ACB211CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"ACB211DCB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"ACB141ABB000", 
x"ACB221CAB000", 
x"ACBD2211CABD", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CBD141CAD000", 
x"ACB141ADB000", 
x"CBD141CAD000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"ACBD2141CCAD", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACBD2111CCBD", 
x"C1C000000000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"ACBD2141CCCD", 
x"CBD141CCD000", 
x"B1B000000000", 
x"CBD141CCD000", 
x"ACBD2141CCDD", 
x"C1C000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"ACB211DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"B1B000000000", 
x"CBD141CDD000", 
x"CBD141CDD000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"ACB141ABB000", 
x"ACB221DAB000", 
x"ACBD2211DABD", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AC21DC000000", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"ACBD2141DCAD", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACBD2111DCBD", 
x"AC21DC000000", 
x"ACB211CCB000", 
x"AC21DC000000", 
x"ACBD2141DCCD", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACBD2141DCDD", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACCA1221AAAA", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACCA1241AABA", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"ACCA1211AACA", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"ACCA1241AADA", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"ACCA1421ABAA", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACCA1411ABCA", 
x"ACC141ABC000", 
x"CC11CC000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"ACCA1121ACAA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCA1141ACBA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCA1111ACCA", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACCA1141ACDA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCA1421ADAA", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACCA1411ADCA", 
x"ACC141ADC000", 
x"ACC211DCC000", 
x"ACC141ADC000", 
x"ACCA1441ADDA", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"AC11AC000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"ACCA2111CCCA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"AC11AC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"ACCA2141DCBA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACCA2111DCCA", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACCA2141DCDA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"ACCB1221AAAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"CCB221AAB000", 
x"ACCB1241AABB", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"AC11AC000000", 
x"ACCB1211AACB", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACCB1241AADB", 
x"ACC141ADC000", 
x"A1A000000000", 
x"CB21AB000000", 
x"ACCB1421ABAB", 
x"AC11AC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"ACCB1411ABCB", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"ACCB1121ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CCB211ACB000", 
x"ACCB1141ACBB", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"ACC111ACC000", 
x"ACCB1111ACCB", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"ACCB1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACCB1421ADAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"ACCB1411ADCB", 
x"ACC211DCC000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"ACCB1441ADDB", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"CCB211ACB000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CCB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"ACC211DCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACCB2221CAAB", 
x"AC11AC000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"AC11AC000000", 
x"ACCB2211CACB", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"ACCB2121CCAB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"ACCB2111CCCB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC3B1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACCB2221DAAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"ACCB2211DACB", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACCB2121DCAB", 
x"AC11AC000000", 
x"AC21DC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"ACC211DCC000", 
x"ACCB2111DCCB", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"ACCB2141DCDB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"CB11CB000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"ACC141ABC000", 
x"ACCC1411ABCC", 
x"ACC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCC1121ACAC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCC1141ACBC", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACCC1111ACCC", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCC1141ACDC", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"ACC141ADC000", 
x"ACCC1411ADCC", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACCC1441ADDC", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACC141ABC000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCC121CAC000", 
x"ACC111ACC000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACC141ADC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCC141CBC000", 
x"CC11CC000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"CCC141CDC000", 
x"ACC211DCC000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACCC2121DCAC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACCC2141DCBC", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACCC2111DCCC", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACCC2141DCDC", 
x"AC21DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"000000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACCD1221AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"ACCD1241AABD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"ACCD1211AACD", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"ACCD1241AADD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACCD1421ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"ACC141ABC000", 
x"CC11CC000000", 
x"ACCD1411ABCD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCD1121ACAD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCD1141ACBD", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACCD1111ACCD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACCD1141ACDD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACCD1421ADAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"ACC141ADC000", 
x"ACC211DCC000", 
x"ACCD1411ADCD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"ACCD1441ADDD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACC141ABC000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"ACCD2111CCCD", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"ACC211DCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC11AC000000", 
x"ACCD2121DCAD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACCD2141DCBD", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACCD2111DCCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACDA1221AAAA", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"ACDA1241AABA", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACDA1211AADA", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACDA1421ABAA", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACDA1441ABBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"ACDA1411ABDA", 
x"ACD141ABD000", 
x"AC21DC000000", 
x"ACD141ABD000", 
x"ACDA1121ACAA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDA1141ACBA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDA1141ACCA", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDA1111ACDA", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"AC11AC000000", 
x"CDA211ADA000", 
x"ACDA1441ADBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"ACDA1411ADDA", 
x"ACD141ADD000", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"CDA211ADA000", 
x"A1A000000000", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"AC11AC000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACDA2211CADA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"AC11AC000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDA2121CCAA", 
x"CDA141CCA000", 
x"AC11AC000000", 
x"CDA141CCA000", 
x"ACDA2141CCBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDA2141CCCA", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"ACDA2111CCDA", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACDA2121DCAA", 
x"AC21DC000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ACDA2141DCBA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACDA2141DCCA", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211CCD000", 
x"ACDA2111DCDA", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ACDB1221AAAB", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"CDB221AAB000", 
x"ACDB1241AABB", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"AC11AC000000", 
x"ACDB1141AC3B", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD121AAD000", 
x"ACDB1211AADB", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"DB21AB000000", 
x"ACDB1421ABAB", 
x"AC11AC000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ACDB1441ABBB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"ACDB1411ABDB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"ACDB1121ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDB1141AC3B", 
x"ACDB1141ACBB", 
x"ACDB1141AC3B", 
x"ACDB1141AC3B", 
x"AC11AC000000", 
x"ACDB1141ACCB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACDB1111ACDB", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"ACDB1421ADAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"AC21DC000000", 
x"ACDB1441ADCB", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"ACD141ADD000", 
x"ACDB1411ADDB", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACDB1141AC3B", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CCB000", 
x"B1B000000000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACD211DCD000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACDB2221CAAB", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"AC11AC000000", 
x"ACDB1141AC3B", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"C1C000000000", 
x"ACDB2211CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACDB2121CCAB", 
x"AC11AC000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"ACDB2141CCBB", 
x"CDB141CCB000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"ACDB2141CCCB", 
x"C1C000000000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACDB2111CCDB", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD3B1141CDAB", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD3B1141CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"ACDB2221DAAB", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"ACDB1141AC3B", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"ACDB2211DADB", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"ACDB2121DCAB", 
x"AC11AC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"ACDB2141DCBB", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACDB2141DCCB", 
x"AC21DC000000", 
x"ACD211CCD000", 
x"ACD211DCD000", 
x"ACDB2111DCDB", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACDC1241AABC", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACDC1211AADC", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACDC1441ABBC", 
x"A1A000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"ACD141ABD000", 
x"ACD141ABD000", 
x"ACDC1411ABDC", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDC1121ACAC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDC1141ACBC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDC1141ACCC", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACDC1111ACDC", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACDC1441ADBC", 
x"A1A000000000", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"ACD211DCD000", 
x"ACD141ADD000", 
x"ACD141ADD000", 
x"ACDC1411ADDC", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"CDC211ADC000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"ACD111ACD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDC2211CADC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDC2121CCAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDC2141CCBC", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACDC2111CCDC", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACDC2211DADC", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ACDC2121DCAC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ACDC2141DCBC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ACDC2141DCCC", 
x"ACD211CCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACDC2111DCDC", 
x"ACD211DCD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACDD1241AABD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACDD1211AADD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACDD1421ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACDD1441ABBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"ACD141ABD000", 
x"ACD141ABD000", 
x"AC21DC000000", 
x"ACDD1411ABDD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDD1121ACAD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDD1141ACBD", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACDD1141ACCD", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACDD1111ACDD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACDD1421ADAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACDD1441ADBD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"ACDD1411ADDD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"CDD211ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"ACDD2121CCAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACDD2141CCBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACDD2111CCDD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC21DC000000", 
x"ACDD2211DADD", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"DD11DD000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC11AC000000", 
x"ACDD2121DCAD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACDD2141DCBD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACD211CCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACDD2111DCDD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AC11AC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ACD211DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADAA1211AAAA", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAA1411ABAA", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"AD11AD000000", 
x"ADAA1441ABBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAA1421ABCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAA1411ACAA", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"AD11AD000000", 
x"ADAA1441ACBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAA1421ACCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA211CDA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAA1111ADAA", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADAA1141ADBA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAA1121ADCA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAA1121ADDA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADA121AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADAA2111CDAA", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"AD11AD000000", 
x"ADAA2141CDBA", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADAA2121CDCA", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211DDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211CDA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADAA2111DDAA", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"AD11AD000000", 
x"ADAA2141DDBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADAA2121DDCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"ADAB1211AAAB", 
x"ADA121AAA000", 
x"AD11AD000000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"ADA141ACA000", 
x"ADAB1221AACB", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"ADAB1221AADB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AB11AB000000", 
x"ADAB1411ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ADA141ACA000", 
x"ADAB1411ACAB", 
x"ADA141ACA000", 
x"AD11AD000000", 
x"DAB221ACB000", 
x"ADAB1441ACBB", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"ADAB1421ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA211CDA000", 
x"ADAB1421ACDB", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"ADAB1111ADAB", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADAB1141AD3B", 
x"ADAB1141ADBB", 
x"ADAB1141AD3B", 
x"ADAB1141AD3B", 
x"AD11AD000000", 
x"ADAB1121ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAB1121ADDB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADA111ADA000", 
x"ADAB1141AD3B", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADA121AAA000", 
x"ADAB2211CAAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ADA141ACA000", 
x"ADAB2221CACB", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"ADAB1141AD3B", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"AB21DB000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"ADAB2111CDAB", 
x"ADA211CDA000", 
x"AD11AD000000", 
x"AB21DB000000", 
x"ADAB2141CDBB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"ADAB2121CDCB", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211DDA000", 
x"ADAB2121CDDB", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"ADAB2211DAAB", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA3B1141DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADA111ADA000", 
x"ADAB1141AD3B", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211CDA000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"ADAB2111DDAB", 
x"ADA211DDA000", 
x"AD11AD000000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"A1A000000000", 
x"ADAB2121DDCB", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"ADAB2121DDDB", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"ADAC1211AAAC", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"ADAC1241AABC", 
x"A1A000000000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"ADAC1221AADC", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"ADAC1411ABAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAC1441ABBC", 
x"A1A000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADAC1421ABCC", 
x"C1C000000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"ADAC1421ABDC", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ADAC1411ACAC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADAC1111ADAC", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAC1141ADBC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAC1121ADCC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAC1121ADDC", 
x"AD11AD000000", 
x"ADA121AAA000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA211CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"AC21DC000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"C1C000000000", 
x"ADAC2211CAAC", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA211CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"ADAC2111CDAC", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADAC2141CDBC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADAC2121CDCC", 
x"C1C000000000", 
x"ADA211DDA000", 
x"C1C000000000", 
x"ADAC2121CDDC", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADAC2211DAAC", 
x"AD11AD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC11AC000000", 
x"AD11AD000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"ADA211CDA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"ADAC2111DDAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADAC2141DDBC", 
x"D1D000000000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"ADAC2121DDDC", 
x"D1D000000000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"ADAD1211AAAD", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1241AABD", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1221AACD", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"ADAD1411ABAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1441ABBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1421ABCD", 
x"DA11DA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1421ABDD", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"ADAD1411ACAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1441ACBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1421ACCD", 
x"ADA211CDA000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADAD1421ACDD", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADAD1111ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAD1141ADBD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAD1121ADCD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADAD1121ADDD", 
x"ADA121AAA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DDD000", 
x"ADA121AAA000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"ADAD2111CDAD", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADAD2141CDBD", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADAD2121CDCD", 
x"ADA211DDA000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADAD2121CDDD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADA111ADA000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211CDA000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"ADAD2111DDAD", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADAD2141DDBD", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADAD2121DDCD", 
x"ADA211DDA000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"ADBA1241AAAA", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADBA1211AABA", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADBA1241AACA", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"ADBA1411ABBA", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADBA1441ACAA", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADBA1411ACBA", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADBA1441ACDA", 
x"ADB211CDB000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADBA1141ADAA", 
x"AD3B1141ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADBA1111ADBA", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADBA1141ADCA", 
x"AD3B1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADBA1141ADDA", 
x"ADB211DDB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB121AAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ADB111ADB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADBA2211CABA", 
x"ADB141ABB000", 
x"ADB221CAB000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADBA2141CDAA", 
x"ADB221DAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADBA2111CDBA", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADBA2141CDCA", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADBA2141CDDA", 
x"ADB211DDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DBA141DAA000", 
x"ADB121AAB000", 
x"DBA141DAA000", 
x"AD11AD000000", 
x"ADBA2211DABA", 
x"ADB141ABB000", 
x"ADB221DAB000", 
x"ADB221DAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"ADB221CAB000", 
x"DBA141DCA000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"ADB221DAB000", 
x"DBA141DDA000", 
x"AD11AD000000", 
x"ADBA2111DDBA", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADBA2141DDCA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADBA2141DDDA", 
x"ADB211DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB121AAB000", 
x"ADBB1211AABB", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB21AB000000", 
x"DB3B2141ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"ADBB1411ABBB", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB3B2141ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"ADBB1441ACAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB141ACB000", 
x"ADBB1411ACBB", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADBB1141ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADBB1111ADBB", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"ADBB1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADBB1141ADDB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"DBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBB141DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DBB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB221CAB000", 
x"ADBB2211CABB", 
x"ADB221CAB000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADBB2141CDAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB211CDB000", 
x"ADBB2111CDBB", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"ADBB2141CDCB", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DBB141DAB000", 
x"ADBB2211DABB", 
x"DBB141DAB000", 
x"DBB141DAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"DB3B1141DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB3B1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB3B1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DBB141DCB000", 
x"BB11BB000000", 
x"DBB141DCB000", 
x"DBB141DCB000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADBB2141DDAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"ADBB2111DDBB", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"A1A000000000", 
x"ADBB2141DDCB", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"ADBC1241AAAC", 
x"AD11AD000000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADBC1211AABC", 
x"ADB121AAB000", 
x"C1C000000000", 
x"ADB141ACB000", 
x"ADBC1241AACC", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADBC1241AADC", 
x"AD11AD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADBC1411ABBC", 
x"ADB141ABB000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"ADB221CAB000", 
x"ADBC1441ACAC", 
x"AD11AD000000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADBC1411ACBC", 
x"ADB141ACB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADB211CDB000", 
x"ADBC1441ACDC", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD3B1141ADAB", 
x"ADBC1141ADAC", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADBC1111ADBC", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD3B1141ADCB", 
x"ADBC1141ADCC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"ADBC1141ADDC", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ABB000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ADB121AAB000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB221CAB000", 
x"ADB141ABB000", 
x"ADBC2211CABC", 
x"ADB221CAB000", 
x"C1C000000000", 
x"ADB141ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ADB221CAB000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADB211CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADB221DAB000", 
x"ADBC2141CDAC", 
x"AD11AD000000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADBC2111CDBC", 
x"ADB211CDB000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADBC2141CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"ADB211DDB000", 
x"ADBC2141CDDC", 
x"C1C000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB221DAB000", 
x"ADB141ABB000", 
x"ADBC2211DABC", 
x"ADB221DAB000", 
x"DBC141DAC000", 
x"ADB141ACB000", 
x"DBC141DAC000", 
x"DBC141DAC000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"ADB221CAB000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"ADB211CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ADB221DAB000", 
x"ADBC2141DDAC", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADBC2111DDBC", 
x"ADB211DDB000", 
x"DBC141DDC000", 
x"B1B000000000", 
x"DBC141DDC000", 
x"DBC141DDC000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"ADBC2141DDDC", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADBD1211AABD", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"ADBD1241AACD", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADBD1411ABBD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DB11DB000000", 
x"DBD211ABD000", 
x"DBD211ABD000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADBD1411ACBD", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"ADBD1441ACDD", 
x"AD11AD000000", 
x"AD3B1141ADAB", 
x"AD11AD000000", 
x"ADBD1141ADAD", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADBD1111ADBD", 
x"AD11AD000000", 
x"AD3B1141ADCB", 
x"AD11AD000000", 
x"ADBD1141ADCD", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"AD11AD000000", 
x"ADBD1141ADDD", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"B1B000000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"ADB211DDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB221CAB000", 
x"ADB141ABB000", 
x"ADB221CAB000", 
x"ADBD2211CABD", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB221DAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADBD2111CDBD", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"ADBD2141CDCD", 
x"A1A000000000", 
x"ADB211DDB000", 
x"AD21CD000000", 
x"ADBD2141CDDD", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB221DAB000", 
x"ADB141ABB000", 
x"ADB221DAB000", 
x"ADBD2211DABD", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"ADB211CDB000", 
x"DBD141DCD000", 
x"DBD141DCD000", 
x"A1A000000000", 
x"ADB221DAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADBD2111DDBD", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"ADBD2141DDCD", 
x"DBD141DDD000", 
x"ADB211DDB000", 
x"DBD141DDD000", 
x"DBD141DDD000", 
x"ADCA1221AAAA", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"ADCA1241AABA", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"ADCA1211AACA", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"ADCA1421ABAA", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"ADCA1441ABBA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ADCA1411ABCA", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADCA1441ABDA", 
x"A1A000000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADCA1411ACCA", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC211CDC000", 
x"DC21AC000000", 
x"ADCA1121ADAA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCA1141ADBA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCA1111ADCA", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADCA1141ADDA", 
x"AD11AD000000", 
x"ADC211DDC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"A1A000000000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ADC121AAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ADC111ADC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"ADCA2121CDAA", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADCA2111CDCA", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211DDC000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"ADCA2211DACA", 
x"ADC221DAC000", 
x"ADC141ACC000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"DCA141DBA000", 
x"DCA141DBA000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ADCA2121DDAA", 
x"DCA141DDA000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"ADCA2141DDBA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ADCA2111DDCA", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADCA2141DDDA", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADCB1221AAAB", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"DCB221AAB000", 
x"ADCB1241AABB", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"ADC121AAC000", 
x"ADCB1211AACB", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"ADCB1241AADB", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"CB21AB000000", 
x"ADCB1421ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"ADCB1441ABBB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"ADCB1411ABCB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"ADCB1441ABDB", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"ADCB1421ACAB", 
x"DC21AC000000", 
x"AD11AD000000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"ADC141ACC000", 
x"ADCB1411ACCB", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"DC21AC000000", 
x"ADCB1441ACDB", 
x"ADC211CDC000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"ADCB1121ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCB1141AD3B", 
x"ADCB1141ADBB", 
x"ADCB1141AD3B", 
x"ADCB1141AD3B", 
x"ADC111ADC000", 
x"ADCB1111ADCB", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"ADCB1141ADDB", 
x"ADC211DDC000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADCB1141AD3B", 
x"ADC111ADC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"ADC211DDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"ADCB2221CAAB", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"ADCB2211CACB", 
x"ADC141ACC000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADCB1141AD3B", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADCB2121CDAB", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADCB2141CDBB", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"ADCB2111CDCB", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"ADCB2141CDDB", 
x"ADC211DDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"ADCB2221DAAB", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"ADC221DAC000", 
x"ADCB2211DACB", 
x"ADC141ACC000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"ADCB1141AD3B", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC3B1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"ADCB2121DDAB", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"ADC211DDC000", 
x"ADCB2111DDCB", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"A1A000000000", 
x"ADCB2141DDDB", 
x"ADC211DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADCC1211AACC", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADCC1421ABAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADCC1441ABBC", 
x"A1A000000000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADCC1411ABCC", 
x"ADC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADCC1421ACAC", 
x"AD11AD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"ADCC1411ACCC", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC211CDC000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCC1121ADAC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCC1141ADBC", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADCC1111ADCC", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCC1141ADDC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DCC121DAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC141ABC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADCC2211CACC", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADCC2121CDAC", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADCC2141CDBC", 
x"C1C000000000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADCC2111CDCC", 
x"ADC211CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211DDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"DCC121DAC000", 
x"DCC121DAC000", 
x"ADCC2211DACC", 
x"DCC121DAC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"DCC141DBC000", 
x"CC11CC000000", 
x"DCC141DBC000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADCC2121DDAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADCC2141DDBC", 
x"D1D000000000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADCC2111DDCC", 
x"ADC211DDC000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"ADCD1241AABD", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADCD1211AACD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ADCD1441ABBD", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADCD1411ABCD", 
x"A1A000000000", 
x"A1A000000000", 
x"DC11DC000000", 
x"ADCD1441ABDD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADCD1411ACCD", 
x"DCD211ACD000", 
x"DCD211ACD000", 
x"ADC211CDC000", 
x"DCD211ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCD1121ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADCD1141ADBD", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADCD1111ADCD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC211DDC000", 
x"ADCD1141ADDD", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"DCD211ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"ADC211CDC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"DCD141DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC141ABC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC141ACC000", 
x"ADCD2211CACD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"ADC211CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADCD2111CDCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"ADC211DDC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"ADC221DAC000", 
x"ADC221DAC000", 
x"ADC141ACC000", 
x"ADCD2211DACD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCD141DBD000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"ADCD2141DDBD", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADCD2111DDCD", 
x"DCD141DDD000", 
x"DCD141DDD000", 
x"ADC211DDC000", 
x"DCD141DDD000", 
x"ADDA1221AAAA", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADDA1241AABA", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"ADDA1241AACA", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"ADDA1211AADA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADDA1421ABAA", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADDA1441ABBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDA1441ABCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDA1411ABDA", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"DD11DD000000", 
x"ADDA1421ACAA", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADDA1441ACBA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDA1441ACCA", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDA1411ACDA", 
x"ADD141ACD000", 
x"ADD141ACD000", 
x"ADD211CDD000", 
x"ADDA1121ADAA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDA1141ADBA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDA1141ADCA", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDA1111ADDA", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA141DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"ADDA2141CDBA", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADDA2141CDCA", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADDA2111CDDA", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADD211CDD000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADDA2111DDDA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"ADDB1221AAAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"DDB221AAB000", 
x"ADDB1241AABB", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"A1A000000000", 
x"ADDB1241AACB", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"ADDB1211AADB", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"DB21AB000000", 
x"ADDB1421ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADDB1441ABBB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADDB1441ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADDB1411ABDB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"ADDB1421ACAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADDB1441ACBB", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADDB1441ACCB", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"ADDB1411ACDB", 
x"ADD141ACD000", 
x"ADD211CDD000", 
x"AD11AD000000", 
x"ADDB1121ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DDB211ADB000", 
x"ADDB1141ADBB", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"AD11AD000000", 
x"ADDB1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADDB1111ADDB", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"ADD111ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADDB2221CAAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"ADDB2211CADB", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"ADDB2121CDAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"A1A000000000", 
x"ADDB2141CDCB", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"ADDB2111CDDB", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"ADDB2221DAAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"ADDB2211DADB", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"ADD211CDD000", 
x"DD11DD000000", 
x"ADDB2121DDAB", 
x"DD11DD000000", 
x"AD11AD000000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"ADDB2141DDCB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADDB2111DDDB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDC1221AAAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDC1241AABC", 
x"ADD141ABD000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"ADDC1241AACC", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDC1211AADC", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDC1421ABAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDC1441ABBC", 
x"A1A000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADDC1441ABCC", 
x"C1C000000000", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"ADDC1411ABDC", 
x"DD11DD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADDC1421ACAC", 
x"AD11AD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADDC1441ACBC", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADDC1441ACCC", 
x"DC21AC000000", 
x"ADD141ACD000", 
x"ADD141ACD000", 
x"ADDC1411ACDC", 
x"ADD211CDD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDC1121ADAC", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDC1141ADBC", 
x"AD11AD000000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"ADDC1141ADCC", 
x"DDC211ADC000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADDC1111ADDC", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DDC221AAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DDC211ADC000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DDC121DAC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDC2211CADC", 
x"ADD111ADD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"ADD211CDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADDC2121CDAC", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADDC2141CDBC", 
x"C1C000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADDC2111CDDC", 
x"ADD211CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDC2221DAAC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDC2211DADC", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADDC2121DDAC", 
x"AD11AD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADDC2141DDBC", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"ADDC2111DDDC", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDD1441ABBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDD1441ABCD", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"ADDD1411ABDD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDD1441ACBD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADDD1441ACCD", 
x"ADD141ACD000", 
x"ADD141ACD000", 
x"ADD141ACD000", 
x"ADDD1411ACDD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDD1121ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDD1141ADBD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADDD1141ADCD", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADDD1111ADDD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADDD2141CDBD", 
x"A1A000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADDD2141CDCD", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"ADDD2111CDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DDD141DCD000", 
x"DDD141DCD000", 
x"ADD211CDD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AD11AD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAAA1111BAAA", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAAA1141BABA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAA1121BACA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAA1121BADA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1211BCAA", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1221BCCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1221BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1211BDAA", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1221BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAA1221BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAA111AAA000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAA121ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AAA111AAA000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAA121ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAA121ADA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AAB121ACB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB121ADB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BAA111BAA000", 
x"BAAB1411B3AB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAA121BCA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAA121BDA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAAB1111BAAB", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAAB1411B3AB", 
x"BAAB1141BABB", 
x"BAAB1411B3AB", 
x"BAAB1411B3AB", 
x"BA11BA000000", 
x"BAAB1121BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAB1121BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"BAAB1411BBAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAB1441BBBB", 
x"BAAB1441B3BB", 
x"BAAB1441B3BB", 
x"BAA121BCA000", 
x"BAAB1421BBCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAAB1421BBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAAB1211BCAB", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BA11BA000000", 
x"BAAB1241BCBB", 
x"BAAB1421B3CB", 
x"BAAB1421B3CB", 
x"B1B000000000", 
x"BAAB1221BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAB1221BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAAB1211BDAB", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BA11BA000000", 
x"BAAB1241BDBB", 
x"BAAB1421B3DB", 
x"BAAB1421B3DB", 
x"B1B000000000", 
x"BAAB1221BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAB1221BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAAB1411B3AB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAB1441B3BB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAAB1421B3CB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAAB1421B3DB", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAAB1411B3AB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAB1441B3BB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAAB1421B3CB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAAB1421B3DB", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC121ADC000", 
x"AA11AA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC121ADC000", 
x"B1B000000000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAAC1111BAAC", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAC1141BABC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAC1121BACC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAC1121BADC", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BAAC1411BBAC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAAC1441BBBC", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"BAAC1421BBCC", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"BAAC1421BBDC", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAAC1211BCAC", 
x"BAA121BCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAAC1241BCBC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAC1221BCCC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAC1221BCDC", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAAC1211BDAC", 
x"BAA121BDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAAC1241BDBC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAC1221BDCC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAC1221BDDC", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC211CAC000", 
x"B1B000000000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"AAC121ADC000", 
x"C1C000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC211CAC000", 
x"AC21DC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"AAC221DDC000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAC221DDC000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"B1B000000000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAAD1111BAAD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAD1141BABD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAD1121BACD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAD1121BADD", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAAD1411BBAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1441BBBD", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1421BBCD", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1421BBDD", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAAD1211BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1241BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1221BCCD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1221BCDD", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAAD1211BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1241BDBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1221BDCD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAAD1221BDDD", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211CAD000", 
x"B1B000000000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AAD221CCD000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAD221CCD000", 
x"AAD221CCD000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD211DAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"AAD211DAD000", 
x"B1B000000000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AAD211DAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"ABA141AAA000", 
x"ABA141AAA000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"BAB111BAB000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"BABA1411B3BA", 
x"BAB141BBB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAB121BCB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAB121BDB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABA141ACA000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"AB11AB000000", 
x"ABA141ADA000", 
x"ABA141ADA000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BABA1141BAAA", 
x"B3AB1411BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABA1111BABA", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BABA1141BACA", 
x"BA3B1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABA1141BADA", 
x"BA3B1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABA1411B3BA", 
x"BAB111BAB000", 
x"BABA1411B3BA", 
x"BABA1411B3BA", 
x"BABA1411BBBA", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB121BCB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB121BDB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BABA1241BCAA", 
x"B3AB1411BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BABA1211BCBA", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BABA1241BCCA", 
x"B3AB1421BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BABA1241BCDA", 
x"B3AB1421BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BABA1241BDAA", 
x"B3AB1411BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BABA1211BDBA", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BABA1241BDCA", 
x"B3AB1421BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BABA1241BDDA", 
x"B3AB1421BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABA1411B3BA", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"ABA141AAA000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABA141ADA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABA1411B3BA", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"BAB121BCB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAB121BDB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"ABB141ACB000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"ABB141ADB000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BABB1141BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BABB1111BABB", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BABB1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BABB1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"BAB111BAB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BABB1411B3BB", 
x"BABB1411BBBB", 
x"BABB1411B3BB", 
x"BABB1411B3BB", 
x"BB11BB000000", 
x"BAB121BCB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BAB121BDB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BABB1241BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"BABB1211BCBB", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"BABB1241BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BABB1241BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BABB1241BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"BABB1211BDBB", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"BABB1241BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BABB1241BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"BABB1411B3BB", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"BABB1411B3BB", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ABB211DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"B1B000000000", 
x"ABC141AAC000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BABC1411B3BC", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"BAB121BCB000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"BAB121BDB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211CBC000", 
x"B1B000000000", 
x"ABC141ACC000", 
x"B1B000000000", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"ABC141ADC000", 
x"B1B000000000", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3AB1411BAAB", 
x"BABC1141BAAC", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BABC1111BABC", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA3B1141BACB", 
x"BABC1141BACC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA3B1141BADB", 
x"BABC1141BADC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BABC1441BBAC", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BABC1411BBBC", 
x"BAB141BBB000", 
x"BABC1411B3BC", 
x"BAB121BCB000", 
x"BABC1411B3BC", 
x"BABC1411B3BC", 
x"BAB141B3B000", 
x"BAB121BDB000", 
x"BABC1441BBDC", 
x"BAB141B3B000", 
x"BC11BC000000", 
x"B3AB1411BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BABC1211BCBC", 
x"BAB121BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3AB1411BDAB", 
x"BABC1241BDAC", 
x"B1B000000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BABC1211BDBC", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B3AB1421BDCB", 
x"BABC1241BDCC", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1421BDDB", 
x"BABC1241BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"C1C000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ABC141ADC000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BABC1411B3BC", 
x"BAB141B3B000", 
x"ABC211CBC000", 
x"BAB121BCB000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211CBC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BABC1411B3BC", 
x"BAB141B3B000", 
x"ABC211DBC000", 
x"BAB121BCB000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211CBC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"ABD141AAD000", 
x"B1B000000000", 
x"ABD141AAD000", 
x"ABD141AAD000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"AB11AB000000", 
x"BABD1411B3BD", 
x"AB11AB000000", 
x"BAB121BCB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"BAB121BDB000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"B1B000000000", 
x"ABD141ACD000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"B1B000000000", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"BA11BA000000", 
x"B3AB1411BAAB", 
x"BA11BA000000", 
x"BABD1141BAAD", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BABD1111BABD", 
x"BA11BA000000", 
x"BA3B1141BACB", 
x"BA11BA000000", 
x"BABD1141BACD", 
x"BA11BA000000", 
x"BA3B1141BADB", 
x"BA11BA000000", 
x"BABD1141BADD", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BABD1411BBBD", 
x"BAB141B3B000", 
x"BAB121BCB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BABD1411B3BD", 
x"BAB121BDB000", 
x"BABD1411B3BD", 
x"BABD1411B3BD", 
x"B1B000000000", 
x"B3AB1411BCAB", 
x"B1B000000000", 
x"BABD1241BCAD", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BABD1211BCBD", 
x"B1B000000000", 
x"B3AB1421BCCB", 
x"B1B000000000", 
x"BABD1241BCCD", 
x"B1B000000000", 
x"B3AB1421BCDB", 
x"B1B000000000", 
x"BABD1241BCDD", 
x"BD11BD000000", 
x"B3AB1411BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BABD1211BDBD", 
x"BD11BD000000", 
x"B3AB1421BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3AB1421BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BABD1411B3BD", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"BAB121BDB000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ABD141ADD000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BABD1411B3BD", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211DBD000", 
x"BAB121BDB000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"ABD211DBD000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ACA121AAA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACA121AAA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA111ACA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BACA1411B3CA", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211DCA000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BACA1121BAAA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACA1141BABA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACA1111BACA", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BACA1141BADA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BACA1411BBCA", 
x"BAC141BBC000", 
x"BAC121BCC000", 
x"BAC141BBC000", 
x"BACA1441BBDA", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"BACA1411B3CA", 
x"BACA1411B3CA", 
x"B3AC1411BCAC", 
x"BACA1411B3CA", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACA1211BCCA", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BACA1241BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACA1221BDAA", 
x"B1B000000000", 
x"B3AC1411BDAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACA1211BDCA", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BACA1241BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA111ACA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BACA1411B3CA", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"ACA211CCA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACA211CCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211CCA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211DCA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA121AAA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA111ACA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BACA1411B3CA", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"ACA211DCA000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACA211DCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211CCA000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACA211DCA000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BACB1141BA3B", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACB1441BB3B", 
x"BAC141BBC000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"BACB1411B3CB", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACB1241BD3B", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC3B1141ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"ACB211CCB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BACB1121BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACB1141BA3B", 
x"BACB1141BABB", 
x"BACB1141BA3B", 
x"BACB1141BA3B", 
x"BAC111BAC000", 
x"BACB1111BACB", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BACB1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACB1421BBAB", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACB1441BBBB", 
x"BAC141BBC000", 
x"BACB1441BB3B", 
x"BAC141BBC000", 
x"BACB1411BBCB", 
x"BAC121BCC000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BACB1441BBDB", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACB1221BCAB", 
x"B3AC1411BCAC", 
x"B1B000000000", 
x"BACB1411B3CB", 
x"BACB1411B3CB", 
x"BACB1411B3CB", 
x"BACB1411B3CB", 
x"BAC121BCC000", 
x"BACB1211BCCB", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"BACB1241BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACB1221BDAB", 
x"B3AC1411BDAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"BACB1241BDBB", 
x"BACB1241BD3B", 
x"BACB1241BD3B", 
x"BAC121BDC000", 
x"BACB1211BDCB", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"BACB1241BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BACB1141BA3B", 
x"BAC111BAC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BACB1411B3CB", 
x"BAC121BCC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BAC121BDC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB211DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BACB1141BA3B", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACB1441BB3B", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACB1411B3CB", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACB1241BD3B", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"ACB211CCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"B1B000000000", 
x"ACC211DCC000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACC1121BAAC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACC1141BABC", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BACC1111BACC", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACC1141BADC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"BAC141BBC000", 
x"BACC1411BBCC", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACC1221BCAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BACC1241BCBC", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BACC1211BCCC", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACC1241BCDC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACC1221BDAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BACC1241BDBC", 
x"B1B000000000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BACC1211BDCC", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACC1241BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BA11BA000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD121AAD000", 
x"B1B000000000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BACD1411B3CD", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"ACD141ADD000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACD1121BAAD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACD1141BABD", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BACD1111BACD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BACD1141BADD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"BACD1441BBBD", 
x"BAC141BBC000", 
x"BAC141BBC000", 
x"BAC121BCC000", 
x"BACD1411BBCD", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"BACD1441BBDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BCAC", 
x"BACD1221BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACD1241BCBD", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BACD1211BCCD", 
x"BACD1411B3CD", 
x"BACD1411B3CD", 
x"BACD1411B3CD", 
x"BACD1411B3CD", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BDAC", 
x"BACD1221BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACD1241BDBD", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BACD1211BDCD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BACD1241BDDD", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BACD1411B3CD", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"B1B000000000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD121AAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD141ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BACD1411B3CD", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD211CCD000", 
x"ACD211DCD000", 
x"B1B000000000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"B1B000000000", 
x"ADA121AAA000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADA141ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BADA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"ADA141ACA000", 
x"B1B000000000", 
x"ADA141ACA000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA211CDA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BADA1121BAAA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADA1141BABA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADA1141BACA", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADA1111BADA", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"BADA1441BBCA", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BADA1411BBDA", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD121BDD000", 
x"BADA1221BCAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AD1411BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADA1241BCCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADA1211BCDA", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BADA1221BDAA", 
x"BADA1411B3DA", 
x"BADA1411B3DA", 
x"B3AD1411BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADA1241BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADA1211BDDA", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"ADA121AAA000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADA141ACA000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADA111ADA000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BADA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211CDA000", 
x"B1B000000000", 
x"ADA211CDA000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADA211DDA000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADA111ADA000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BADA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211CDA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"B1B000000000", 
x"ADA211DDA000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA211DDA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BADB1141BA3B", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"BADB1241BC3B", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"BADB1411B3DB", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"AD3B1141ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD3B1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BADB1121BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADB1141BA3B", 
x"BADB1141BABB", 
x"BADB1141BA3B", 
x"BADB1141BA3B", 
x"BA11BA000000", 
x"BADB1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BADB1111BADB", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BADB1421BBAB", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BADB1441BBBB", 
x"BADB1441B3BB", 
x"BAD141BBD000", 
x"B1B000000000", 
x"BADB1441BBCB", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"BADB1411BBDB", 
x"BAD141BBD000", 
x"BAD121BDD000", 
x"B1B000000000", 
x"BADB1221BCAB", 
x"B1B000000000", 
x"B3AD1411BCAD", 
x"BA11BA000000", 
x"BADB1241BCBB", 
x"BADB1241BC3B", 
x"BADB1241BC3B", 
x"B1B000000000", 
x"BADB1241BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BADB1211BCDB", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"BADB1221BDAB", 
x"B1B000000000", 
x"B3AD1411BDAD", 
x"BADB1411B3DB", 
x"BADB1241BDBB", 
x"BADB1411B3DB", 
x"BADB1411B3DB", 
x"B1B000000000", 
x"BADB1241BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"BADB1211BDDB", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BADB1141BA3B", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BADB1441B3BB", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"BADB1241BC3B", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"BADB1411B3DB", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BADB1141BA3B", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BAD121BCD000", 
x"DB11DB000000", 
x"BADB1411B3DB", 
x"DB11DB000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB211CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1411B3DC", 
x"BAD121BDD000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC141ACC000", 
x"B1B000000000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"DC21AC000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADC211DDC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADC1121BAAC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADC1141BABC", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADC1141BACC", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BADC1111BADC", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADC1421BBAC", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BADC1441BBBC", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1441BBCC", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BADC1411BBDC", 
x"BAD121BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1221BCAC", 
x"B3AD1411BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"BADC1241BCBC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1241BCCC", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BADC1211BCDC", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1221BDAC", 
x"B3AD1411BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"BADC1241BDBC", 
x"B1B000000000", 
x"BADC1411B3DC", 
x"BADC1411B3DC", 
x"BADC1241BDCC", 
x"BADC1411B3DC", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BADC1211BDDC", 
x"BAD121BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADC141ACC000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1411B3DC", 
x"BAD121BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"B1B000000000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"ADC211DDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ADC121AAC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC221DAC000", 
x"B1B000000000", 
x"ADC141ACC000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADC1411B3DC", 
x"BAD121BDD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ADC221DAC000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADC211DDC000", 
x"B1B000000000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"A1A000000000", 
x"B1B000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"B1B000000000", 
x"ADD141ACD000", 
x"ADD211CDD000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADD1121BAAD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADD1141BABD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BADD1141BACD", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BADD1111BADD", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BADD1411BBDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1221BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1241BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1241BCCD", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BADD1211BCDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1221BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1241BDBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BADD1241BDCD", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BADD1211BDDD", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"ADD211CDD000", 
x"B1B000000000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"ADD211CDD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BAA111BAA000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BAA121BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"B3BA1411BABA", 
x"BB11BB000000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBAA1111BBAA", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAA1121BBCA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAA1121BBDA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAA1411BCAA", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"B3BA1411BCBA", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"BBAA1421BCCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAA1421BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAA1411BDAA", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"B3BA1411BDBA", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"BBAA1421BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAA1421BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BAA121BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BAA121BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBAB1141BB3B", 
x"BB11BB000000", 
x"BB11BB000000", 
x"AB11AB000000", 
x"BAB121BCB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BAB121BDB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BBAB1411BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BBAB1421BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBAB1421BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBAB1111BBAB", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBAB1141BBBB", 
x"BBAB1141BB3B", 
x"BBAB1141BB3B", 
x"BB11BB000000", 
x"BBAB1121BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAB1121BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBAB1411BCAB", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BAB121BCB000", 
x"BB11BB000000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"BBAB1421BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAB1421BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBAB1411BDAB", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BAB121BDB000", 
x"BB11BB000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"BBAB1421BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAB1421BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBAB1141BB3B", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBAB1141BB3B", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBAC1411BAAC", 
x"BA11BA000000", 
x"B3BA1411BABA", 
x"BB11BB000000", 
x"BBAC1441BABC", 
x"B3B141BAB000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBAC1421BADC", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBAC1111BBAC", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BBAC1141BBBC", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAC1121BBCC", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAC1121BBDC", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBAC1411BCAC", 
x"BBA141BCA000", 
x"B3BA1411BCBA", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAC1421BCDC", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBAC1411BDAC", 
x"BBA141BDA000", 
x"B3BA1411BDBA", 
x"BB11BB000000", 
x"BBAC1441BDBC", 
x"B3B141BDB000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAC1421BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBAD1411BAAD", 
x"B3BA1411BABA", 
x"BB11BB000000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBAD1111BBAD", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAD1141BBBD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAD1121BBCD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBAD1121BBDD", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBAD1411BCAD", 
x"B3BA1411BCBA", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAD1421BCCD", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBAD1411BDAD", 
x"B3BA1411BDBA", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBAD1421BDCD", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AD21CD000000", 
x"AD21CD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BBB141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBBA1411BABA", 
x"B3BB1411BABB", 
x"BBB141BAB000", 
x"BBB141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB3B1141BBAB", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBBA1111BBBA", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBBA1141BBCA", 
x"BB3B1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBBA1141BBDA", 
x"BB3B1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3BB1441BCAB", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBBA1411BCBA", 
x"B3BB1411BCBB", 
x"BBB141BCB000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B3BB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBA1441BCDA", 
x"B3BB1441BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"B3BB1441BDAB", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBBA1411BDBA", 
x"B3BB1411BDBB", 
x"BBB141BDB000", 
x"BBB141BDB000", 
x"BBBA1441BDCA", 
x"BB3B1441BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBA1441BDDA", 
x"B3BB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BBB141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BBB141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBBB1441BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"BBBB1411BABB", 
x"BBB141BAB000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BBBB1441BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBB1441BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBBB1141BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBBB1111BBBB", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BBBB1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBBB1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBBB1441BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"BBBB1411BCBB", 
x"BBB141BCB000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"BBBB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBB1441BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBB1441BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"BBBB1411BDBB", 
x"BBB141BDB000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"BBBB1441BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBBB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BBB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3BB1441BAAB", 
x"BBBC1441BAAC", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B3BB1411BABB", 
x"BBBC1411BABC", 
x"BBB141BAB000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"B3BB1441BADB", 
x"BBBC1441BADC", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB3B1141BBAB", 
x"BBBC1141BBAC", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBBC1111BBBC", 
x"BBB111BBB000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BB3B1141BBDB", 
x"BBBC1141BBDC", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BBB141BCB000", 
x"B3BB1411BCBB", 
x"BBBC1411BCBC", 
x"BBB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3BB1441BDAB", 
x"BBBC1441BDAC", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B3BB1411BDBB", 
x"BBBC1411BDBC", 
x"BBB141BDB000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"B3BB1441BDDB", 
x"BBBC1441BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BBB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BBB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BBB141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3BB1441BAAB", 
x"B1B000000000", 
x"BBBD1441BAAD", 
x"BBB141BAB000", 
x"B3BB1411BABB", 
x"BBB141BAB000", 
x"BBBD1411BABD", 
x"B1B000000000", 
x"BB3B1441BACB", 
x"B1B000000000", 
x"BBBD1441BACD", 
x"BBD141BAD000", 
x"B3BB1441BADB", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB3B1141BBAB", 
x"BB11BB000000", 
x"BBBD1141BBAD", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBBD1111BBBD", 
x"BB11BB000000", 
x"BB3B1141BBCB", 
x"BB11BB000000", 
x"BBBD1141BBCD", 
x"BBD111BBD000", 
x"BB3B1141BBDB", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3BB1441BCAB", 
x"B1B000000000", 
x"BBBD1441BCAD", 
x"BBB141BCB000", 
x"B3BB1411BCBB", 
x"BBB141BCB000", 
x"BBBD1411BCBD", 
x"B1B000000000", 
x"B3BB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"B3BB1441BCDB", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BBB141BDB000", 
x"B3BB1411BDBB", 
x"BBB141BDB000", 
x"BBBD1411BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BBB141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BBB141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"B3BC1411BABC", 
x"B3B141BAB000", 
x"BBCA1411BACA", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBCA1441BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCA1121BBAA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCA1141BBBA", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBCA1111BBCA", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBCA1141BBDA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BB11BB000000", 
x"B3BC1411BCBC", 
x"BC11BC000000", 
x"BBCA1411BCCA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BBCA1421BDAA", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3BC1411BDBC", 
x"B3B141BDB000", 
x"BBCA1411BDCA", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBCA1441BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BCA121BAA000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBCB1141BB3B", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBCB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BB11BB000000", 
x"B3BC1411BABC", 
x"BCB121BAB000", 
x"BBC141BAC000", 
x"BBCB1411BACB", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BBCB1441BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBCB1121BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCB1141BB3B", 
x"BBCB1141BBBB", 
x"BBC111BBC000", 
x"BBCB1141BB3B", 
x"BBC111BBC000", 
x"BBCB1111BBCB", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBCB1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BBCB1411BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BBCB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BB11BB000000", 
x"B3BC1411BDBC", 
x"BCB141BDB000", 
x"BBC141BDC000", 
x"BBCB1411BDCB", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"BBCB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BCB121BAB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BB11BB000000", 
x"BBCB1141BB3B", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BCB141BDB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBCB1141BB3B", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCC1421BAAC", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"B3BC1411BABC", 
x"B3B141BAB000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BBCC1411BACC", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCC1441BADC", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCC1121BBAC", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBCC1111BBCC", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCC1141BBDC", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BB11BB000000", 
x"B3BC1411BCBC", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCC1421BDAC", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3BC1411BDBC", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBCC1411BDCC", 
x"BBC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCC1441BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"BCD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCD1421BAAD", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"B3BC1411BABC", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBCD1411BACD", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCD1121BBAD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BBCD1141BBBD", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBCD1111BBCD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBCD1141BBDD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BB11BB000000", 
x"B3BC1411BCBC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BBCD1411BCCD", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBCD1421BDAD", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3BC1411BDBC", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBCD1411BDCD", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"BCD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"BCD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BDA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BDA111BDA000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"B3B141BAB000", 
x"B3BD1411BABD", 
x"BBDA1441BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDA1411BADA", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BBDA1121BBAA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDA1141BBBA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBDA1141BBCA", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDA1111BBDA", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3BD1411BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDA1411BCDA", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3BD1411BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BBDA1411BDDA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BDA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BDA111BDA000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"BDA121BAA000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BDA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BDA111BDA000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBDB1141BB3B", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BB11BB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BBDB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BB11BB000000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BBDB1441BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BBDB1411BADB", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBDB1121BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDB1141BB3B", 
x"BBDB1141BBBB", 
x"BBDB1141BB3B", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BBDB1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBDB1111BBDB", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BBDB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"BB11BB000000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"BBDB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BBDB1411BCDB", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BBDB1421BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BBDB1441BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BBDB1411BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BBDB1141BB3B", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BB11BB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BDB121BAB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BB11BB000000", 
x"BBDB1141BB3B", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"DB11DB000000", 
x"BDB141BCB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BB11BB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BDC121BAC000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BDC141BCC000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDC1421BAAC", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"BBDC1441BABC", 
x"B3BD1411BABD", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BBDC1411BADC", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDC1121BBAC", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDC1141BBBC", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDC1141BBCC", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBDC1111BBDC", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDC1421BCAC", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3BD1411BCBD", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BBDC1411BCDC", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BBDC1421BDAC", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"BBDC1441BDBC", 
x"B3BD1411BDBD", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BBDC1411BDDC", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BDC121BAC000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BDC141BCC000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BDC121BAC000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BDC141BCC000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDD1421BAAD", 
x"B3B141BAB000", 
x"BB11BB000000", 
x"B3B141BAB000", 
x"B3BD1411BABD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDD1441BACD", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BBDD1411BADD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDD1121BBAD", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBDD1141BBCD", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBDD1111BBDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBDD1421BCAD", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3BD1411BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BBDD1411BCDD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3BD1411BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCAA1211BAAA", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCAA1241BABA", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CA1411BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAA1221BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAA1411BBAA", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAA1111BCAA", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCAA1141BCBA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAA1121BCCA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAA1121BCDA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAA1411BDAA", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCAA1441BDBA", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CA1411BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAA1421BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"BC11BC000000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCAB1411B3AB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"BCA111BCA000", 
x"BCAB1141BC3B", 
x"BC11BC000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCAB1211BAAB", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCAB1411B3AB", 
x"BCAB1241BABB", 
x"BCAB1411B3AB", 
x"BCAB1411B3AB", 
x"B3CA1411BACA", 
x"BCAB1221BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAB1221BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA121BAA000", 
x"BCAB1411BBAB", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCAB1441B3BB", 
x"BCAB1441BBBB", 
x"BC11BC000000", 
x"BCAB1441B3BB", 
x"BCA111BCA000", 
x"BCAB1141BC3B", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCAB1421BBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCAB1111BCAB", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCAB1141BC3B", 
x"BCAB1141BCBB", 
x"BCAB1141BC3B", 
x"BCAB1141BC3B", 
x"BC11BC000000", 
x"BCAB1121BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAB1121BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCAB1411BDAB", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCAB1421B3DB", 
x"BCAB1441BDBB", 
x"BC11BC000000", 
x"BCAB1421B3DB", 
x"B3CA1411BDCA", 
x"BCAB1421BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAB1421BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA3B1141CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA3B1141CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BCA121BAA000", 
x"BCAB1411B3AB", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"BC11BC000000", 
x"CAB141CBB000", 
x"BCA111BCA000", 
x"BCAB1141BC3B", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCAB1421B3DB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"BC11BC000000", 
x"CAB121CCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"BC11BC000000", 
x"CAB121CDB000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCAB1411B3AB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"BCAB1441B3BB", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCAB1141BC3B", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCAB1421B3DB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"BCAC1411B3AC", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC121CCC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCAC1211BAAC", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CA1411BACA", 
x"BCAC1411B3AC", 
x"BCAC1221BACC", 
x"BCAC1411B3AC", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAC1221BADC", 
x"B1B000000000", 
x"BCA121BAA000", 
x"BCA141BBA000", 
x"BCAC1411BBAC", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"BCAC1421BBDC", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCAC1111BCAC", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAC1141BCBC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAC1121BCCC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAC1121BCDC", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCAC1411BDAC", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CA1411BDCA", 
x"B1B000000000", 
x"BCAC1421BDCC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAC1421BDDC", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"BCAC1411B3AC", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"BCAC1411B3AC", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"B1B000000000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1411B3AD", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCAD1211BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCAD1241BABD", 
x"B3CA1411BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1221BACD", 
x"BCAD1411B3AD", 
x"BCAD1411B3AD", 
x"BCAD1411B3AD", 
x"BCAD1221BADD", 
x"BCA121BAA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCAD1411BBAD", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCAD1441BBBD", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1421BBDD", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCAD1111BCAD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAD1141BCBD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAD1121BCCD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCAD1121BCDD", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCAD1411BDAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCAD1441BDBD", 
x"B3CA1411BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1421BDCD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1421BDDD", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1411B3AD", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"B1B000000000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"B1B000000000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCAD1411B3AD", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"BCB121BAB000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"BCBA1411B3BA", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3CB1421BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BCBA1211BABA", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BA11BA000000", 
x"B3CB1411BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BC3B1241BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BCBA1411B3BA", 
x"BCB121BAB000", 
x"BCBA1411B3BA", 
x"BCBA1411B3BA", 
x"BCBA1411BBBA", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BCB141BDB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCBA1141BCAA", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCBA1111BCBA", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCBA1141BCCA", 
x"B3CB1411BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCBA1141BCDA", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCBA1441BDAA", 
x"B3CB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCBA1411BDBA", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCBA1441BDDA", 
x"B3CB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CBA141CAA000", 
x"CBA211ABA000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"BCB121BAB000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"BCBA1411B3BA", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BCB141BDB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CAA000", 
x"B1B000000000", 
x"CBA141CCA000", 
x"CBA141CCA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"CBA141CDA000", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BCB121BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BCBA1411B3BA", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBB211ABB000", 
x"BCBB1411B3BB", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCBB1241BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BCBB1211BABB", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCBB1241BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BCB121BAB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BCBB1411B3BB", 
x"BCBB1411BBBB", 
x"BCBB1411B3BB", 
x"BCBB1411B3BB", 
x"BB11BB000000", 
x"BCB111BCB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BCBB1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCBB1111BCBB", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BCBB1141BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCBB1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCBB1441BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BCBB1411BDBB", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCBB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BCB121BAB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BCBB1411B3BB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCBC1411B3BC", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3CB1421BAAB", 
x"BCBC1241BAAC", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCBC1211BABC", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"BCBC1241BACC", 
x"B1B000000000", 
x"B1B000000000", 
x"BC3B1241BADB", 
x"BCBC1241BADC", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB121BAB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCBC1411BBBC", 
x"BCB141BBB000", 
x"BCBC1411B3BC", 
x"BCB111BCB000", 
x"BCBC1411B3BC", 
x"BCBC1411B3BC", 
x"BCB141B3B000", 
x"BCB141BDB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BCBC1141BCAC", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCBC1111BCBC", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"B3CB1411BCCB", 
x"BCBC1141BCCC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BCBC1141BCDC", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CB1421BDAB", 
x"BCBC1441BDAC", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCBC1411BDBC", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"BCBC1441BDCC", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CB1441BDDB", 
x"BCBC1441BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CAC000", 
x"CB11CB000000", 
x"CBC141CAC000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BCB121BAB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BCB141BBB000", 
x"BCBC1411B3BC", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"BCB111BCB000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BCB141BDB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CB11CB000000", 
x"CBC141CDC000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCBC1411B3BC", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCBD1411B3BD", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CBD211ABD000", 
x"BCB141BDB000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3CB1421BAAB", 
x"B1B000000000", 
x"BCBD1241BAAD", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCBD1211BABD", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"B1B000000000", 
x"BCBD1241BACD", 
x"B1B000000000", 
x"BC3B1241BADB", 
x"B1B000000000", 
x"BCBD1241BADD", 
x"BCB141B3B000", 
x"BCB121BAB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCBD1411BBBD", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCBD1411B3BD", 
x"BCB141BDB000", 
x"BCBD1411B3BD", 
x"BCBD1411B3BD", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BCBD1141BCAD", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCBD1111BCBD", 
x"BC11BC000000", 
x"B3CB1411BCCB", 
x"BC11BC000000", 
x"BCBD1141BCCD", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BCBD1141BCDD", 
x"BD11BD000000", 
x"B3CB1421BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCBD1411BDBD", 
x"BD11BD000000", 
x"B3CB1411BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"B1B000000000", 
x"CBD141CAD000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"BCB121BAB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCBD1411B3BD", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"CBD141CCD000", 
x"B1B000000000", 
x"CBD141CCD000", 
x"CBD141CDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"B1B000000000", 
x"CBD141CDD000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCBD1411B3BD", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"BCB141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCA211ACA000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CCA211ACA000", 
x"B1B000000000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCCA1221BAAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCA1241BABA", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCA1211BACA", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCCA1241BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCA1421BBAA", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCA1411BBCA", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BCCA1121BCAA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCA1141BCBA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCA1111BCCA", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCCA1141BCDA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCA1421BDAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCA1411BDCA", 
x"BCC141BDC000", 
x"B3CC1411BDCC", 
x"BCC141BDC000", 
x"BCCA1441BDDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BC11BC000000", 
x"CC11CC000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"B1B000000000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCA211ACA000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCCB1421B3AB", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCB1441B3BB", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCCB1411B3CB", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCB1441B3DB", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"BC11BC000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCCB1221BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCB1421B3AB", 
x"BCCB1241BABB", 
x"BC11BC000000", 
x"BCCB1421B3AB", 
x"BCC121BAC000", 
x"BCCB1211BACB", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"BCCB1241BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCB1421BBAB", 
x"BCC121BAC000", 
x"B1B000000000", 
x"BCCB1441B3BB", 
x"BCCB1441BBBB", 
x"BC11BC000000", 
x"BCCB1441B3BB", 
x"BC11BC000000", 
x"BCCB1411BBCB", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCB1441BBDB", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCCB1121BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCB1411B3CB", 
x"BCCB1141BCBB", 
x"BCCB1411B3CB", 
x"BCCB1411B3CB", 
x"BCC111BCC000", 
x"BCCB1111BCCB", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BCCB1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCB1441B3DB", 
x"BCCB1441BDBB", 
x"BC11BC000000", 
x"BCCB1441B3DB", 
x"BCC141BDC000", 
x"BCCB1411BDCB", 
x"B3CC1411BDCC", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BCCB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"BC11BC000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BCC121BAC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BCCB1411B3CB", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB121CAB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC3B1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"BC11BC000000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCCB1421B3AB", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCB1441B3BB", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCCB1411B3CB", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCCB1441B3DB", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCC1221BAAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCCC1211BACC", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCC1241BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCC1121BCAC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCC1141BCBC", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCCC1111BCCC", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCC1141BCDC", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCC1421BDAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"BCC141BDC000", 
x"BCCC1411BDCC", 
x"BCC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCC1441BDDC", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCC121CAC000", 
x"CCC121CAC000", 
x"CC11CC000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BC11BC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CCC141CDC000", 
x"CCC141CDC000", 
x"CC11CC000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD221AAD000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD211ACD000", 
x"B1B000000000", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCD1221BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCCD1241BABD", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCCD1211BACD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCD1241BADD", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"BCCD1421BBAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BCCD1411BBCD", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCD1121BCAD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCD1141BCBD", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCCD1111BCCD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCCD1141BCDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCD1421BDAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"BCC141BDC000", 
x"B3CC1411BDCC", 
x"BCCD1411BDCD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCCD1441BDDD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BC11BC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCDA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"CDA121CAA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDA141CCA000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"B1B000000000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"BCDA1221BAAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDA1241BABA", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCDA1241BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCDA1211BADA", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCDA1421BBAA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"BCDA1441BBBA", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCDA1411BBDA", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BDD000", 
x"BCDA1121BCAA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDA1141BCBA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDA1141BCCA", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDA1111BCDA", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCDA1421BDAA", 
x"BCDA1411B3DA", 
x"BCDA1411B3DA", 
x"BCDA1411B3DA", 
x"BCDA1441BDBA", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCDA1441BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCDA1411BDDA", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"CDA121CAA000", 
x"B1B000000000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCDA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"CDA121CAA000", 
x"B1B000000000", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDA141CCA000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCDA1411B3DA", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"CDA121CAA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDA141CCA000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"BCDB1421B3AB", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"BCDB1441B3BB", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BCDB1141BC3B", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"BCDB1411B3DB", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"BC11BC000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"BCDB1221BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDB1421B3AB", 
x"BCDB1241BABB", 
x"BC11BC000000", 
x"BCDB1421B3AB", 
x"B1B000000000", 
x"BCDB1241BACB", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"BCDB1211BADB", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"BCDB1421BBAB", 
x"B1B000000000", 
x"BCD121BAD000", 
x"BCDB1441B3BB", 
x"BCDB1441BBBB", 
x"BC11BC000000", 
x"BCDB1441B3BB", 
x"BC11BC000000", 
x"BCDB1141BC3B", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"BCDB1411BBDB", 
x"BCD141BBD000", 
x"BCD141BDD000", 
x"BC11BC000000", 
x"BCDB1121BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDB1141BC3B", 
x"BCDB1141BCBB", 
x"BCDB1141BC3B", 
x"BCDB1141BC3B", 
x"BC11BC000000", 
x"BCDB1141BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCDB1111BCDB", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"BCDB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDB1411B3DB", 
x"BCDB1411B3DB", 
x"BCDB1411B3DB", 
x"BCDB1411B3DB", 
x"B1B000000000", 
x"BCDB1441BDCB", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"BCDB1411BDDB", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"BC11BC000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCDB1421B3AB", 
x"B1B000000000", 
x"BCD121BAD000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"BCDB1141BC3B", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"BCDB1411B3DB", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD3B1141CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD3B1141CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BCD121BAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"BCDB1141BC3B", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"DB11DB000000", 
x"BCDB1411B3DB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1411B3DC", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1221BAAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1241BACC", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCDC1211BADC", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1421BBAC", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCDC1411BBDC", 
x"BCD141BDD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDC1121BCAC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDC1141BCBC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDC1141BCCC", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCDC1111BCDC", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1421BDAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCDC1411B3DC", 
x"BCDC1411B3DC", 
x"BCDC1411B3DC", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCDC1411BDDC", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1411B3DC", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDC1411B3DC", 
x"BCD141BDD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"CDC121CAC000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD211ADD000", 
x"B1B000000000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDD1221BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCDD1241BABD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCDD1211BADD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCDD1411BBDD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDD1121BCAD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDD1141BCBD", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCDD1141BCCD", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCDD1111BCDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCDD1421BDAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCDD1441BDBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCDD1411BDDD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAA121DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDAA1211BAAA", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDAA1241BABA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDAA1221BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAA1221BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAA1411BBAA", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDAA1421BBCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAA1411BCAA", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDAA1441BCBA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDAA1421BCCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAA1421BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAA1111BDAA", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDAA1141BDBA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAA1121BDCA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAA1121BDDA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAA121DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DAA121DCA000", 
x"B1B000000000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAA121DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDAB1411B3AB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BDA111BDA000", 
x"BDAB1141BD3B", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDAB1211BAAB", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDAB1411B3AB", 
x"BDAB1241BABB", 
x"BDAB1411B3AB", 
x"BDAB1411B3AB", 
x"B1B000000000", 
x"BDAB1221BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BADA", 
x"BDAB1221BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA121BAA000", 
x"BDAB1411BBAB", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDAB1441BBBB", 
x"BDAB1441B3BB", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDAB1421BBCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDAB1421BBDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDAB1411BCAB", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDAB1421B3CB", 
x"BDAB1441BCBB", 
x"BDAB1421B3CB", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDAB1421BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BCDA", 
x"BDAB1421BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDAB1111BDAB", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDAB1141BD3B", 
x"BDAB1141BDBB", 
x"BDAB1141BD3B", 
x"BDAB1141BD3B", 
x"BD11BD000000", 
x"BDAB1121BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAB1121BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDAB1411B3AB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"BDAB1441B3BB", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDAB1421B3CB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDAB1141BD3B", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB211AAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA3B1141DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA3B1141DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"BDA121BAA000", 
x"BDAB1411B3AB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDAB1421B3CB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDAB1141BD3B", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"DAC211AAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAC211AAC000", 
x"B1B000000000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC221ADC000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"BDAC1411B3AC", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAC221ADC000", 
x"B1B000000000", 
x"DAC121DCC000", 
x"DAC221ADC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDAC1211BAAC", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAC1241BABC", 
x"BD11BD000000", 
x"BDAC1411B3AC", 
x"BDAC1411B3AC", 
x"BDAC1221BACC", 
x"BDAC1411B3AC", 
x"B3DA1411BADA", 
x"B1B000000000", 
x"BDAC1221BADC", 
x"B1B000000000", 
x"BDA121BAA000", 
x"BDA141BBA000", 
x"BDAC1411BBAC", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"BDAC1441BBBC", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"BDAC1421BBCC", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BDAC1421BBDC", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDAC1411BCAC", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAC1441BCBC", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAC1421BCCC", 
x"B1B000000000", 
x"B3DA1411BCDA", 
x"B1B000000000", 
x"BDAC1421BCDC", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDAC1111BDAC", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAC1141BDBC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAC1121BDCC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAC1121BDDC", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DAC211AAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"BDAC1411B3AC", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DAC121DCC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"BDAC1411B3AC", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAC121DCC000", 
x"B1B000000000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAC121DDC000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1411B3AD", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDAD1211BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1221BACD", 
x"B3DA1411BADA", 
x"BDAD1411B3AD", 
x"BDAD1411B3AD", 
x"BDAD1221BADD", 
x"BDA121BAA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDAD1411BBAD", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1421BBCD", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDAD1411BCAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1421BCCD", 
x"B3DA1411BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1421BCDD", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDAD1111BDAD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAD1141BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAD1121BDCD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDAD1121BDDD", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1411B3AD", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DAD121DDD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDAD1411B3AD", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"BDB121BAB000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"BDBA1411B3BA", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B3DB1421BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BDBA1211BABA", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BA11BA000000", 
x"BD3B1241BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B3DB1411BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BDBA1411B3BA", 
x"BDB121BAB000", 
x"BDBA1411B3BA", 
x"BDBA1411B3BA", 
x"BDBA1411BBBA", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDB141BCB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDBA1441BCAA", 
x"B3DB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDBA1411BCBA", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B3DB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDBA1441BCDA", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDBA1141BDAA", 
x"BD3B1141BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDBA1111BDBA", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDBA1141BDCA", 
x"BD3B1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDBA1141BDDA", 
x"B3DB1411BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BDB121BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BDBA1411B3BA", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"B1B000000000", 
x"DBA141DAA000", 
x"DBA141DAA000", 
x"DBA211ABA000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"BDB121BAB000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"BDBA1411B3BA", 
x"BDB141BBB000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BDB141BCB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"DBA141DCA000", 
x"DBA141DCA000", 
x"BA11BA000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"B1B000000000", 
x"DBA141DDA000", 
x"DBA141DDA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DBB211ABB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBB211ABB000", 
x"BDBB1411B3BB", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDBB1241BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BDBB1211BABB", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BDBB1241BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDBB1241BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BDB121BAB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BDBB1411B3BB", 
x"BDBB1411BBBB", 
x"BDBB1411B3BB", 
x"BDBB1411B3BB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BDB111BDB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BDBB1441BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"BDBB1411BCBB", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"BDBB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDBB1141BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDBB1111BDBB", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BDBB1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDBB1141BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DBB211ABB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BDBB1411B3BB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"DBB211ABB000", 
x"DBB141DAB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BDB121BAB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"BDB141BCB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"BB11BB000000", 
x"DBB141DCB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"DBC211ABC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDBC1411B3BC", 
x"BD11BD000000", 
x"DBC211ABC000", 
x"BDB141BCB000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3DB1421BAAB", 
x"BDBC1241BAAC", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDBC1211BABC", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BD3B1241BACB", 
x"BDBC1241BACC", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BADB", 
x"BDBC1241BADC", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB121BAB000", 
x"BDBC1441BBAC", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDBC1411BBBC", 
x"BDB141BBB000", 
x"BDBC1411B3BC", 
x"BDBC1411B3BC", 
x"BDBC1411B3BC", 
x"BDBC1411B3BC", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDBC1441BBDC", 
x"BD11BD000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDBC1411BCBC", 
x"BDB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B3DB1411BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"BD3B1141BDAB", 
x"BDBC1141BDAC", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDBC1111BDBC", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD3B1141BDCB", 
x"BDBC1141BDCC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3DB1411BDDB", 
x"BDBC1141BDDC", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"DBC211ABC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDBC1411B3BC", 
x"BD11BD000000", 
x"BC11BC000000", 
x"BDB141BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"DBC211ABC000", 
x"BD11BD000000", 
x"DBC141DAC000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BDB121BAB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BDB141BBB000", 
x"BDBC1411B3BC", 
x"BD11BD000000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BC11BC000000", 
x"BD11BD000000", 
x"DBC141DCC000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"BD11BD000000", 
x"DBC141DDC000", 
x"B1B000000000", 
x"DBC141DDC000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDBD1411B3BD", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"B1B000000000", 
x"B3DB1421BAAB", 
x"B1B000000000", 
x"BDBD1241BAAD", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDBD1211BABD", 
x"B1B000000000", 
x"BD3B1241BACB", 
x"B1B000000000", 
x"BDBD1241BACD", 
x"B1B000000000", 
x"B3DB1411BADB", 
x"B1B000000000", 
x"BDBD1241BADD", 
x"BDB141B3B000", 
x"BDB121BAB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDBD1411BBBD", 
x"BDB141B3B000", 
x"BDB141BCB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BDBD1411B3BD", 
x"BDB111BDB000", 
x"BDBD1411B3BD", 
x"BDBD1411B3BD", 
x"B1B000000000", 
x"B3DB1421BCAB", 
x"B1B000000000", 
x"BDBD1441BCAD", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDBD1411BCBD", 
x"B1B000000000", 
x"B3DB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"BDBD1441BCDD", 
x"BD11BD000000", 
x"BD3B1141BDAB", 
x"BD11BD000000", 
x"BDBD1141BDAD", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDBD1111BDBD", 
x"BD11BD000000", 
x"BD3B1141BDCB", 
x"BD11BD000000", 
x"BDBD1141BDCD", 
x"BD11BD000000", 
x"B3DB1411BDDB", 
x"BD11BD000000", 
x"BDBD1141BDDD", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDBD1411B3BD", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBD141DAD000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"BDB121BAB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BDB141BBB000", 
x"DB11DB000000", 
x"BDBD1411B3BD", 
x"DB11DB000000", 
x"BDB141BCB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BDB111BDB000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DB11DB000000", 
x"DBD141DCD000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DBD141DDD000", 
x"DB11DB000000", 
x"DBD141DDD000", 
x"DBD141DDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCA211ACA000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDCA1411B3CA", 
x"B1B000000000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DCA211ACA000", 
x"B1B000000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"DCA121DAA000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCA111DCA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"BDCA1221BAAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCA1241BABA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDCA1211BACA", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDCA1241BADA", 
x"B1B000000000", 
x"B3DC1411BADC", 
x"B1B000000000", 
x"BDCA1421BBAA", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"BDCA1441BBBA", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDCA1411BBCA", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BDCA1411B3CA", 
x"BDCA1411B3CA", 
x"BDCA1411B3CA", 
x"BDCA1411B3CA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDCA1411BCCA", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDCA1441BCDA", 
x"B1B000000000", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BDCA1121BDAA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCA1141BDBA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCA1111BDCA", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDCA1141BDDA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDCA1411B3CA", 
x"B1B000000000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCA111DCA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"B1B000000000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCA211ACA000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDCA1411B3CA", 
x"B1B000000000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA121DAA000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCA141DDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCA111DCA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDCB1421B3AB", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCB1441BB3B", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDCB1411B3CB", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDCB1141BD3B", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"CB11CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDCB1221BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCB1421B3AB", 
x"BDCB1241BABB", 
x"BDCB1421B3AB", 
x"BD11BD000000", 
x"BDC121BAC000", 
x"BDCB1211BACB", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"BDCB1241BADB", 
x"B3DC1411BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCB1421BBAB", 
x"BDC121BAC000", 
x"B1B000000000", 
x"BDCB1441BB3B", 
x"BDCB1441BBBB", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"BDCB1411BBCB", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDCB1441BBDB", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDCB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCB1411B3CB", 
x"BDCB1411B3CB", 
x"BDCB1411B3CB", 
x"BDCB1411B3CB", 
x"BDC141BCC000", 
x"BDCB1411BCCB", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BDCB1441BCDB", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDCB1121BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCB1141BD3B", 
x"BDCB1141BDBB", 
x"BDCB1141BD3B", 
x"BDCB1141BD3B", 
x"BDC111BDC000", 
x"BDCB1111BDCB", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BDCB1141BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BDC121BAC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BDCB1411B3CB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BDCB1141BD3B", 
x"BDC111BDC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDCB1421B3AB", 
x"BDC121BAC000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"BDCB1441BB3B", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDCB1411B3CB", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDCB1141BD3B", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC3B1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1411B3CC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1221BAAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1241BABC", 
x"BD11BD000000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDCC1211BACC", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1241BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDCC1411BBCC", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1421BCAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1441BCBC", 
x"BD11BD000000", 
x"BDCC1411B3CC", 
x"BDCC1411B3CC", 
x"BDCC1411BCCC", 
x"BDCC1411B3CC", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCC1121BDAC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCC1141BDBC", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDCC1111BDCC", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCC1141BDDC", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCC211ACC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1411B3CC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BD11BD000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCC121DAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCC121DAC000", 
x"B1B000000000", 
x"DCC211ACC000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCC1411B3CC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BCC000", 
x"BDCD1411B3CD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"CD11CD000000", 
x"DCD211ACD000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCD1221BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDCD1211BACD", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BADC", 
x"BDCD1241BADD", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"BDCD1421BBAD", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDCD1411BBCD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDCD1421BCAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDCD1411BCCD", 
x"BDCD1411B3CD", 
x"BDCD1411B3CD", 
x"B3DC1411BCDC", 
x"BDCD1411B3CD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCD1121BDAD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCD1141BDBD", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDCD1111BDCD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDCD1141BDDD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DCD211ACD000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BCC000", 
x"BDCD1411B3CD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"DCD121DAD000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD121DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BCC000", 
x"BDCD1411B3CD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD141DDD000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA211ADA000", 
x"B1B000000000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"BDDA1221BAAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDA1241BABA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDDA1241BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDA1211BADA", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDDA1421BBAA", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDDA1441BBBA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDDA1441BBCA", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDDA1411BBDA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDDA1421BCAA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDA1441BCBA", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDDA1441BCCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDA1411BCDA", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDDA1121BDAA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDA1141BDBA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDA1141BDCA", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDA1111BDDA", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"DDA141DCA000", 
x"B1B000000000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"BDDB1421B3AB", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"BDDB1441B3BB", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDDB1441B3CB", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BDDB1411B3DB", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"BDDB1221BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDB1421B3AB", 
x"BDDB1241BABB", 
x"BDDB1421B3AB", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDDB1241BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDDB1211BADB", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"BDDB1421BBAB", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDDB1441B3BB", 
x"BDDB1441BBBB", 
x"BDDB1441B3BB", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDDB1441BBCB", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BDDB1411BBDB", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"B1B000000000", 
x"BDDB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDB1441B3CB", 
x"BDDB1441BCBB", 
x"BDDB1441B3CB", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDDB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDDB1411BCDB", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BDDB1121BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDB1411B3DB", 
x"BDDB1141BDBB", 
x"BDDB1411B3DB", 
x"BDDB1411B3DB", 
x"BD11BD000000", 
x"BDDB1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDDB1111BDDB", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"BDDB1421B3AB", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"BDDB1441B3BB", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDDB1441B3CB", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BDDB1411B3DB", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BDD121BAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDDB1411B3DB", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB121DAB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDB141DCB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"B1B000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDC221AAC000", 
x"B1B000000000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDC211ADC000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1221BAAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1241BABC", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1241BACC", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDDC1211BADC", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1421BBAC", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1441BBBC", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1441BBCC", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDC1411BBDC", 
x"BDD111BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1421BCAC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1441BCBC", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDC1441BCCC", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDDC1411BCDC", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDC1121BDAC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDC1141BDBC", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDC1141BDCC", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDDC1111BDDC", 
x"BDD111BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DDC121DAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDC121DAC000", 
x"B1B000000000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DDC121DAC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDD1221BAAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDD1241BACD", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDDD1211BADD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDD1421BCAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDDD1441BCCD", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDDD1411BCDD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDD1121BDAD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDD1141BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDDD1141BDCD", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDDD1111BDDD", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"B1B000000000", 
x"DDD121DAD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"B1B000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CA11CA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAAA1111CAAA", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAAA1141CABA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAA1121CACA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAA1121CADA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAA1411CBAA", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAAA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAA1421CBDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAA1211CDAA", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAAA1241CDBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAA1221CDDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAA121ADA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AA11AA000000", 
x"CAAB2111AAAB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"CA11CA000000", 
x"CAAB2121AACB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CAAB2121AADB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CAA111CAA000", 
x"CAAB2211ACAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"CA11CA000000", 
x"CAAB2221ACCB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAAB2221ACDB", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"CAAB2211ADAB", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"CA11CA000000", 
x"CAAB2221ADCB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAAB2221ADDB", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"AAB211CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA121CDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAA111CAA000", 
x"CAAB1111CAAB", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"AAB211CAB000", 
x"CAAB1141CABB", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"CA11CA000000", 
x"CAAB1121CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAB1121CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CAAB1411CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAAB1441CBBB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAAB1421CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAAB1421CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAA111CAA000", 
x"CAAB1211CCAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAB221CCB000", 
x"CAAB1241CCBB", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"CA11CA000000", 
x"CAAB1221CCCB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAAB1221CCDB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAAB1211CDAB", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"AAB221CDB000", 
x"CAAB1241CDBB", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"CA11CA000000", 
x"CAAB1221CDCB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAB1221CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"CA11CA000000", 
x"AAB121ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB121ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CAA111CAA000", 
x"AAB211CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"CA11CA000000", 
x"AAB221CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"AAB221CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AAB211DAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"CA11CA000000", 
x"AAB221DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AAB221DDB000", 
x"C1C000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CAAC2111AAAC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CAAC2141AABC", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CAAC2121AADC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAA121CDA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"CAAC2211ADAC", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAAC1111CAAC", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAC1141CABC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAC1121CACC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAC1121CADC", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAAC1411CBAC", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAC1441CBBC", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAAC1421CBCC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAC1421CBDC", 
x"C1C000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CAAC1211CCAC", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"CAAC1241CCBC", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAAC1221CCCC", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"CAAC1221CCDC", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAAC1211CDAC", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAC1241CDBC", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAAC1221CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAC1221CDDC", 
x"C1C000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC121ADC000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AAC211DAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CAAD2111AAAD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CA11CA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AA11AA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CA11CA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AAD141ABD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD121ACD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAAD1111CAAD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAD1141CABD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAD1121CACD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAD1121CADD", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAAD1411CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1441CBBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1421CBCD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1421CBDD", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAAD1211CCAD", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1241CCBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1221CCCD", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1221CCDD", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAAD1211CDAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1241CDBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1221CDCD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAAD1221CDDD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AAD141ABD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAD121ACD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AAD211DAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AAD211DAD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ABA141AAA000", 
x"CAB211AAB000", 
x"ABA141AAA000", 
x"ABA141AAA000", 
x"CABA2111AABA", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABA2141AADA", 
x"CAB221ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CABA2211ACBA", 
x"CAB141CBB000", 
x"CAB221ACB000", 
x"CAB221ACB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABA141ADA000", 
x"AB11AB000000", 
x"ABA141ADA000", 
x"ABA141ADA000", 
x"CABA2211ADBA", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"CAB211AAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ABA211CBA000", 
x"CAB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA211DBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CABA1141CAAA", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CABA1111CABA", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CABA1141CACA", 
x"CA3B1141CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CABA1141CADA", 
x"CA3B1141CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ABA211CBA000", 
x"AB11AB000000", 
x"ABA211CBA000", 
x"ABA211CBA000", 
x"CABA1411CBBA", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CABA1211CCBA", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABA1241CCDA", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABA1241CDAA", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABA1211CDBA", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABA1241CDDA", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABA141AAA000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABA141ADA000", 
x"CAB221ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB11AB000000", 
x"ABA211DBA000", 
x"ABA211DBA000", 
x"BA11BA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ABA211CBA000", 
x"CAB141CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABA211DBA000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"CABB2111AABB", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CABB2141AACB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CABB2141AADB", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB3B1141ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB3B1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB3B1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ABB141ACB000", 
x"CABB2211ACBB", 
x"ABB141ACB000", 
x"ABB141ACB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"CABB2211ADBB", 
x"ABB141ADB000", 
x"ABB141ADB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"ABB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B3B141BCB000", 
x"ABB211CBB000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"ABB211DBB000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CABB1141CAAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CABB1111CABB", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CABB1141CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CABB1141CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CABB1441CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"CABB1411CBBB", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"CA11CA000000", 
x"AB3B2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CABB1441CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CABB1211CCBB", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABB1241CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CABB1211CDBB", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CA11CA000000", 
x"CABB1241CDCB", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CABB1241CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"ABB141ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ABB141ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"CA11CA000000", 
x"AB3B2141DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB3B2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"CABC2141AAAC", 
x"A1A000000000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CABC2111AABC", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"ABC141AAC000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"CABC2141AADC", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"CAB141CBB000", 
x"CABC2211ACBC", 
x"CAB221ACB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CABC2211ADBC", 
x"CAB221ADB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CAB111CAB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CAB121CCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CAB121CDB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB211AAB000", 
x"CABC1141CAAC", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CABC1111CABC", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA3B1141CACB", 
x"CABC1141CACC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA3B1141CADB", 
x"CABC1141CADC", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"CABC1441CBAC", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CABC1411CBBC", 
x"CAB141CBB000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CABC1441CBDC", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CABC1241CCAC", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CABC1211CCBC", 
x"CAB121CCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CABC1241CCCC", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CABC1241CCDC", 
x"C1C000000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"CABC1241CDAC", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CABC1211CDBC", 
x"CAB121CDB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CABC1241CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"CABC1241CDDC", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"ABC141AAC000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"ABC141ADC000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BC11BC000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"CABD2141AAAD", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CABD2111AABD", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABD141AAD000", 
x"CAB221ADB000", 
x"ABD141AAD000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"CAB141CBB000", 
x"CAB221ACB000", 
x"CABD2211ACBD", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CABD2211ADBD", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ABD141ADD000", 
x"AB21DB000000", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"AB11AB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CABD1141CAAD", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CABD1111CABD", 
x"CA11CA000000", 
x"CA3B1141CACB", 
x"CA11CA000000", 
x"CABD1141CACD", 
x"CA11CA000000", 
x"CA3B1141CADB", 
x"CA11CA000000", 
x"CABD1141CADD", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CABD1411CBBD", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CABD1211CCBD", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"CABD1241CCCD", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"CABD1241CCDD", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CABD1241CDAD", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CABD1211CDBD", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CABD1241CDCD", 
x"C1C000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"CABD1241CDDD", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"CA11CA000000", 
x"CAB221ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"C1C000000000", 
x"ABD141ADD000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"BD11BD000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ACA121AAA000", 
x"ACA121AAA000", 
x"CAC211AAC000", 
x"ACA121AAA000", 
x"CACA2141AABA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CACA2111AACA", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"CACA2141AADA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA141ABA000", 
x"ACA141ABA000", 
x"AC11AC000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"CAC111CAC000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAC141CBC000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CAC121CCC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAC121CDC000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"ACA141ADA000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CACA1121CAAA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACA1141CABA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACA1111CACA", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CACA1141CADA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACA1421CBAA", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CACA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACA1411CBCA", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CACA1441CBDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CACA1241CCBA", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CACA1211CCCA", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CACA1241CCDA", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"CACA1221CDAA", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CACA1241CDBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACA1211CDCA", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CACA1241CDDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACA141ADA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CACB2121AAAB", 
x"CAC211AAC000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"CA11CA000000", 
x"CACB2111AACB", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"CACB2141AADB", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB21AB000000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CA11CA000000", 
x"CACB1141CA3B", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"CA11CA000000", 
x"CACB2211ACCB", 
x"CAC121CCC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"CAC121CDC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"CACB2221ADAB", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"CA11CA000000", 
x"CACB2211ADCB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"ACB121AAB000", 
x"CAC211AAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CACB1141CA3B", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CA11CA000000", 
x"ACB211CCB000", 
x"CAC121CCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"ACB211DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CACB1121CAAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACB1141CA3B", 
x"CACB1141CABB", 
x"CACB1141CA3B", 
x"CACB1141CA3B", 
x"CAC111CAC000", 
x"CACB1111CACB", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CACB1141CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CACB1411CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CA11CA000000", 
x"CACB1221CCAB", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"CAC121CCC000", 
x"CACB1211CCCB", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"CACB1241CCDB", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACB1221CDAB", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CACB1241CDBB", 
x"B1B000000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"CACB1211CDCB", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"CACB1241CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB121AAB000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"ACB141ABB000", 
x"ACB221DAB000", 
x"ACB221DAB000", 
x"CA11CA000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CACB1141CA3B", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"CA11CA000000", 
x"ACB211CCB000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"ACB221DAB000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"ACB211DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CACC2141AABC", 
x"A1A000000000", 
x"CA11CA000000", 
x"CAC211AAC000", 
x"CACC2111AACC", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"CACC2141AADC", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"ACC141ABC000", 
x"CC11CC000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAC141CBC000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAC121CDC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"ACC141ADC000", 
x"CACC2211ADCC", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAC121CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACC1121CAAC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACC1141CABC", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CACC1111CACC", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACC1141CADC", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1421CBAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1441CBBC", 
x"C1C000000000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CACC1411CBCC", 
x"CAC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1441CBDC", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAC111CAC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CACC1211CCCC", 
x"CAC121CCC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAC121CDC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1221CDAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1241CDBC", 
x"C1C000000000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CACC1211CDCC", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACC1241CDDC", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ADC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"CAC121CCC000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"CACD2121AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CACD2141AABD", 
x"CA11CA000000", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"CACD2111AACD", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"ACD141ABD000", 
x"ACD141ABD000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CAC141CBC000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CAC121CCC000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACD2211ADCD", 
x"ACD141ADD000", 
x"ACD141ADD000", 
x"C1C000000000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CAC121CDC000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACD1121CAAD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACD1141CABD", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CACD1111CACD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CACD1141CADD", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"CACD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACD1441CBBD", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CACD1411CBCD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CACD1441CBDD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"CACD1241CCBD", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CACD1211CCCD", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CAC121CDC000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CACD1211CDCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"ACD211CCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"CAC121CDC000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211DCD000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"CAD211AAD000", 
x"CADA2141AABA", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADA2111AADA", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CADA2211ACDA", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CA11CA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADA121AAA000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"ADA211CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CADA1121CAAA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADA1141CABA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADA1141CACA", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADA1111CADA", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CADA1421CBAA", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CADA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADA1411CBDA", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CADA1241CCBA", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CADA1211CCDA", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CADA1221CDAA", 
x"ADA211CDA000", 
x"ADA211CDA000", 
x"AD11AD000000", 
x"CADA1241CDBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADA1211CDDA", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CAD211AAD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CA11CA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"ADA211CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"ADA211DDA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADA211DDA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CADB2121AAAB", 
x"C1C000000000", 
x"CAD211AAD000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"CA11CA000000", 
x"CADB2141AACB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"CADB2111AADB", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"CADB1141CA3B", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"CADB2211ACDB", 
x"C1C000000000", 
x"CAD121CDD000", 
x"AD11AD000000", 
x"AD3B1141ADAB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"CA11CA000000", 
x"AD3B1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CADB2211ADDB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CADB1141CA3B", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAD121CCD000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"CAD121CDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CADB1121CAAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADB1141CA3B", 
x"CADB1141CABB", 
x"CADB1141CA3B", 
x"CADB1141CA3B", 
x"CA11CA000000", 
x"CADB1141CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CADB1111CADB", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"CADB1421CBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CADB1441CBBB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CADB1441CBCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CADB1411CBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CADB1221CCAB", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"CADB1241CCBB", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CADB1241CCCB", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CADB1211CCDB", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"CADB1221CDAB", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB211CDB000", 
x"CADB1241CDBB", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"CA11CA000000", 
x"CADB1241CDCB", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"CADB1211CDDB", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"ADB221DAB000", 
x"ADB141ABB000", 
x"ADB221DAB000", 
x"ADB221DAB000", 
x"CA11CA000000", 
x"ADB141ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"CADB1141CA3B", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"ADB211CDB000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"ADB221DAB000", 
x"C1C000000000", 
x"AD11AD000000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"ADB211DDB000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CADC2121AAAC", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"CADC2141AABC", 
x"A1A000000000", 
x"CA11CA000000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CADC2111AADC", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC2211ACDC", 
x"CAD121CDD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CADC2211ADDC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ADC141ACC000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADC1121CAAC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADC1141CABC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADC1141CACC", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CADC1111CADC", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC1421CBAC", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC1441CBBC", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CADC1441CBCC", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CADC1411CBDC", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADC1221CCAC", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC1241CCBC", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CADC1241CCCC", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CADC1211CCDC", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC1221CDAC", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADC1241CDBC", 
x"C1C000000000", 
x"CA11CA000000", 
x"ADC211CDC000", 
x"CADC1241CDCC", 
x"ADC211CDC000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CADC1211CDDC", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"ADC141ACC000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CA11CA000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CAD121CCD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CADD2141AABD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CADD2111AADD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CA11CA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADD1121CAAD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADD1141CABD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CADD1141CACD", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CADD1111CADD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1441CBBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1441CBCD", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CADD1411CBDD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CADD1211CCDD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1221CDAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1241CDBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CADD1241CDCD", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CADD1211CDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ADD141ABD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AD11AD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"CB21AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AA11AA000000", 
x"CB11CB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CBAA2111ABAA", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"BA11BA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAA2121ABCA", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAA2121ABDA", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CB11CB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBAA1411CAAA", 
x"CB21AB000000", 
x"CBA141CAA000", 
x"CBA141CAA000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAA1421CACA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAA1421CADA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAA1111CBAA", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBAA1141CBBA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAA1121CBCA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAA1121CBDA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAA1411CCAA", 
x"CB21AB000000", 
x"CBA141CCA000", 
x"CBA141CCA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAA1411CDAA", 
x"CB21AB000000", 
x"CBA141CDA000", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBAA1421CDCA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAA1421CDDA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"CB21AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CBAB2111ABAB", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"BA11BA000000", 
x"CBAB2141ABBB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CBAB2121ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CBAB2121ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CBA141CAA000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBAB1141CB3B", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3AB1411BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA3B1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA3B1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB121BCB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB121BDB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B3AB1411BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA111CBA000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1421BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1411BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1421BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CBAB1411CAAB", 
x"CBA141CAA000", 
x"CBA141CAA000", 
x"CBA211ABA000", 
x"CBAB1441CABB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAB1421CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBAB1111CBAB", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBAB1141CB3B", 
x"CBAB1141CBBB", 
x"CBAB1141CB3B", 
x"CBAB1141CB3B", 
x"CB11CB000000", 
x"CBAB1121CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAB1121CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CAA000", 
x"CBAB1411CCAB", 
x"CBA141CCA000", 
x"CBA141CCA000", 
x"CBA111CBA000", 
x"CBAB1141CB3B", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"CBAB1421CCDB", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"CBAB1411CDAB", 
x"CBA141CDA000", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"CBAB1441CDBB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBAB1421CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBAB1141CB3B", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB11CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBAC2111ABAC", 
x"CBA211ABA000", 
x"BA11BA000000", 
x"CB21AB000000", 
x"CBAC2141ABBC", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CBAC2121ABCC", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAC2121ABDC", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"AC11AC000000", 
x"CB11CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"CB11CB000000", 
x"BAC121BCC000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BCAC", 
x"B1B000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BAC121BCC000", 
x"CB11CB000000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BDAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"CB11CB000000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"CBAC1411CAAC", 
x"CBA141CAA000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CBAC1441CABC", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB11CB000000", 
x"CBAC1421CACC", 
x"AC11AC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBAC1421CADC", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBAC1111CBAC", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAC1141CBBC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAC1121CBCC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAC1121CBDC", 
x"CB11CB000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"CBAC1411CCAC", 
x"CBA141CCA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"CBAC1421CCCC", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"CBAC1421CCDC", 
x"C1C000000000", 
x"CBA141CDA000", 
x"CB21AB000000", 
x"CBAC1411CDAC", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"CBAC1441CDBC", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBAC1421CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBAC1421CDDC", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB11CB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBAD2111ABAD", 
x"BA11BA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAD2141ABBD", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CBAD2121ABCD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBAD2121ABDD", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CB21AB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"CB11CB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CB11CB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD141BBD000", 
x"BAD121BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AD1411BCAD", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AD1411BDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"CBA141CAA000", 
x"CBAD1411CAAD", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBAD1421CACD", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"CBAD1421CADD", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBAD1111CBAD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAD1141CBBD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAD1121CBCD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBAD1121CBDD", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"CBA141CCA000", 
x"CBAD1411CCAD", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBAD1421CCCD", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBAD1421CCDD", 
x"CBA141CDA000", 
x"CB21AB000000", 
x"CBA141CDA000", 
x"CBAD1411CDAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBAD1421CDCD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBAD1421CDDD", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"CB3B2141ABAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CBBA2111ABBA", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBBA2141ABCA", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBBA2141ABDA", 
x"CB3B2141ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B3BA1411BABA", 
x"CBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"CB11CB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"CBB141CAB000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"B3BA1411BCBA", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"B3BA1411BDBA", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBBA1441CAAA", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1411CABA", 
x"CBB211ABB000", 
x"CBB141CAB000", 
x"CBB141CAB000", 
x"CBBA1441CACA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1441CADA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1141CBAA", 
x"CB3B1141CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBBA1111CBBA", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBBA1141CBCA", 
x"CB3B1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBBA1141CBDA", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBBA1441CCAA", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1411CCBA", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1441CCDA", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1441CDAA", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1411CDBA", 
x"BB11BB000000", 
x"CBB141CDB000", 
x"CBB141CDB000", 
x"CBBA1441CDCA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBA1441CDDA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBBB2141ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CBBB2111ABBB", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CBBB2141ABCB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBBB2141ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3BB1441BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B3BB1411BABB", 
x"BBB141BAB000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3BB1441BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB3B1141BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB3B1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB3B1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CBB141CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"CBB111CBB000", 
x"BBB141BCB000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3BB1441BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B3BB1411BDBB", 
x"BBB141BDB000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3BB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBBB1441CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"CBBB1411CABB", 
x"CBB141CAB000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBB1441CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBBB1141CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBBB1111CBBB", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CBBB1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBBB1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBB1441CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"CBBB1411CDBB", 
x"CBB141CDB000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBBB1441CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB3B2141ABAB", 
x"CBBC2141ABAC", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBBC2111ABBC", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"CB3B2141ABDB", 
x"CBBC2141ABDC", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"CBB211ABB000", 
x"B3BC1411BABC", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"CB11CB000000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"B3BC1411BCBC", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3BC1411BDBC", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"CB11CB000000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBBC1441CAAC", 
x"C1C000000000", 
x"CBB141CAB000", 
x"CBB211ABB000", 
x"CBBC1411CABC", 
x"CBB141CAB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBBC1441CACC", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBBC1441CADC", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB3B1141CBAB", 
x"CBBC1141CBAC", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBBC1111CBBC", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB3B1141CBCB", 
x"CBBC1141CBCC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CBBC1141CBDC", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"CBBC1441CCAC", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBBC1411CCBC", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBBC1441CCCC", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"CBBC1441CCDC", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBBC1441CDAC", 
x"C1C000000000", 
x"CBB141CDB000", 
x"BB11BB000000", 
x"CBBC1411CDBC", 
x"CBB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBBC1441CDCC", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBBC1441CDDC", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB3B2141ABAB", 
x"CB21AB000000", 
x"CBBD2141ABAD", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBBD2111ABBD", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CBBD2141ABCD", 
x"BD11BD000000", 
x"CB3B2141ABDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"CBB211ABB000", 
x"B3B141BAB000", 
x"B3BD1411BABD", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"CBB141CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"B3BD1411BCBD", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"CBB141CDB000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3BD1411BDBD", 
x"BD11BD000000", 
x"CB11CB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBBD1441CAAD", 
x"CBB141CAB000", 
x"CBB211ABB000", 
x"CBB141CAB000", 
x"CBBD1411CABD", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBBD1441CACD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBBD1441CADD", 
x"CB11CB000000", 
x"CB3B1141CBAB", 
x"CB11CB000000", 
x"CBBD1141CBAD", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBBD1111CBBD", 
x"CB11CB000000", 
x"CB3B1141CBCB", 
x"CB11CB000000", 
x"CBBD1141CBCD", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CBBD1141CBDD", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"CBBD1441CCAD", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CBBD1411CCBD", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"CBBD1441CCDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBBD1441CDAD", 
x"CBB141CDB000", 
x"BB11BB000000", 
x"CBB141CDB000", 
x"CBBD1411CDBD", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBBD1441CDCD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBBD1441CDDD", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"B3B141BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBCA2121ABAA", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCA2141ABBA", 
x"CB21AB000000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"CBCA2111ABCA", 
x"CB11CB000000", 
x"CBC211ABC000", 
x"CBC211ABC000", 
x"CBCA2141ABDA", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CA11CA000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"B3CA1411BACA", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA121BAA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CA1411BDCA", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB21AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBCA1411CACA", 
x"CB11CB000000", 
x"CBC141CAC000", 
x"CBC141CAC000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CBCA1121CBAA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCA1141CBBA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCA1111CBCA", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBCA1141CBDA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CA11CA000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBCA1411CCCA", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"CBCA1421CDAA", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBCA1411CDCA", 
x"CB11CB000000", 
x"CBC141CDC000", 
x"CBC141CDC000", 
x"CBCA1441CDDA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBCB2141AB3B", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBCB2121ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCB2141AB3B", 
x"CBCB2141ABBB", 
x"BC11BC000000", 
x"CBCB2141AB3B", 
x"CBC211ABC000", 
x"CBCB2111ABCB", 
x"CBC211ABC000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBCB2141ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBCB1141CB3B", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3CB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC3B1241BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB121BAB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BCB141BDB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"B3CB1411BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CB1441BDDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBCB1421CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBCB2141AB3B", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CBCB1411CACB", 
x"CBC141CAC000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CBCB1441CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBCB1121CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCB1141CB3B", 
x"CBCB1141CBBB", 
x"CBCB1141CB3B", 
x"CBCB1141CB3B", 
x"CBC111CBC000", 
x"CBCB1111CBCB", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBCB1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBCB1421CCAB", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBCB1141CB3B", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CBCB1411CCCB", 
x"CBC141CCC000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"CBCB1441CCDB", 
x"CBC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBCB1421CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CBCB1411CDCB", 
x"CBC141CDC000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"CBCB1441CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBCB2141AB3B", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBCB1141CB3B", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCC2121ABAC", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB11CB000000", 
x"CBCC2111ABCC", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCC2141ABDC", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"CB11CB000000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"CB11CB000000", 
x"B3CC1411BDCC", 
x"BCC141BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBCC1421CAAC", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CB11CB000000", 
x"CBCC1411CACC", 
x"CBC141CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBCC1441CADC", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCC1121CBAC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCC1141CBBC", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBCC1111CBCC", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCC1141CBDC", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB11CB000000", 
x"CBCC1411CCCC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBCC1421CDAC", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CB11CB000000", 
x"CBCC1411CDCC", 
x"CBC141CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBCC1441CDDC", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCD2121ABAD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BC11BC000000", 
x"CBCD2141ABBD", 
x"CBC211ABC000", 
x"CB11CB000000", 
x"CBC211ABC000", 
x"CBCD2111ABCD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBCD2141ABDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BBD000", 
x"BCD141BDD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBCD1421CAAD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CB11CB000000", 
x"CBC141CAC000", 
x"CBCD1411CACD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBCD1441CADD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCD1121CBAD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCD1141CBBD", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBCD1111CBCD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBCD1141CBDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"CBCD1421CCAD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CBCD1411CCCD", 
x"CD11CD000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CB21AB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CB11CB000000", 
x"CBC141CDC000", 
x"CBCD1411CDCD", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CBDA2121ABAA", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDA2141ABBA", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"CBDA2141ABCA", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDA2111ABDA", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"DA11DA000000", 
x"CB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BADA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA121BAA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BCDA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CB11CB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CBDA1421CAAA", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBDA1441CACA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBDA1411CADA", 
x"B1B000000000", 
x"CBD141CAD000", 
x"CBD141CAD000", 
x"CBDA1121CBAA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDA1141CBBA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDA1141CBCA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDA1111CBDA", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBDA1421CCAA", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"CBDA1411CCDA", 
x"B1B000000000", 
x"CBD141CCD000", 
x"CBD141CDD000", 
x"CBDA1421CDAA", 
x"CB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"CBDA1441CDCA", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBDA1411CDDA", 
x"B1B000000000", 
x"CBD141CDD000", 
x"CBD141CDD000", 
x"DA11DA000000", 
x"CB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"DA11DA000000", 
x"CB11CB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"DA11DA000000", 
x"CB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CBDB2141AB3B", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CBDB2121ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDB2141AB3B", 
x"CBDB2141ABBB", 
x"CBDB2141AB3B", 
x"BD11BD000000", 
x"CB21AB000000", 
x"CBDB2141ABCB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBDB2111ABDB", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CBDB1141CB3B", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3DB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB121BAB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDB141BCB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B3DB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"CBDB1141CB3B", 
x"BDB141BCB000", 
x"CBD111CBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD3B1141BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD3B1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3DB1411BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CBDB1421CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBDB1441CABB", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CBDB1411CADB", 
x"CBD141CAD000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CBDB1121CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDB1141CB3B", 
x"CBDB1141CBBB", 
x"CBDB1141CB3B", 
x"CBDB1141CB3B", 
x"CB11CB000000", 
x"CBDB1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CBDB1111CBDB", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CBDB1421CCAB", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CBDB1141CB3B", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"CBD141CCD000", 
x"CBDB1411CCDB", 
x"CBD141CCD000", 
x"CBD141CDD000", 
x"C1C000000000", 
x"CBDB1421CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"CBDB1441CDBB", 
x"DB11DB000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"CBDB1411CDDB", 
x"CBD141CDD000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CBDB2141AB3B", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"BDB121BAB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BDB141BBB000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BDB141BCB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CBDB1141CB3B", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDC2121ABAC", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDC2141ABBC", 
x"BD11BD000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CBDC2141ABCC", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBDC2111ABDC", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"BDC121BAC000", 
x"CB11CB000000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"CB11CB000000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"BDC141BCC000", 
x"CB11CB000000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBDC1421CAAC", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDC1441CABC", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBDC1441CACC", 
x"C1C000000000", 
x"CBD141CAD000", 
x"B1B000000000", 
x"CBDC1411CADC", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDC1121CBAC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDC1141CBBC", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDC1141CBCC", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBDC1111CBDC", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBDC1421CCAC", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBDC1441CCCC", 
x"CBD141CCD000", 
x"CBD141CCD000", 
x"B1B000000000", 
x"CBDC1411CCDC", 
x"CBD141CDD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBDC1421CDAC", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBDC1441CDBC", 
x"BD11BD000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CBD141CDD000", 
x"B1B000000000", 
x"CBDC1411CDDC", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBDD2121ABAD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CBDD2141ABCD", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBDD2111ABDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CB11CB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBDD1421CAAD", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBDD1441CACD", 
x"CBD141CAD000", 
x"B1B000000000", 
x"CBD141CAD000", 
x"CBDD1411CADD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDD1121CBAD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDD1141CBBD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBDD1141CBCD", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBDD1111CBDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"CBD141CCD000", 
x"B1B000000000", 
x"CBD141CCD000", 
x"CBDD1411CCDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBDD1421CDAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBDD1441CDCD", 
x"CBD141CDD000", 
x"B1B000000000", 
x"CBD141CDD000", 
x"CBDD1411CDDD", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"DD11DD000000", 
x"CB21AB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DD11DD000000", 
x"CB11CB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CCA211ACA000", 
x"AA11AA000000", 
x"CC11CC000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCAA2111ACAA", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCAA2141ACBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAA2121ACDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CC11CC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAA1411CBAA", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CCAA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCAA1421CBDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAA1111CCAA", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCAA1141CCBA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAA1121CCDA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAA1411CDAA", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CCAA1441CDBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCAA1421CDDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"CCAB2211AAAB", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CCA211ACA000", 
x"CCAB2221AACB", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCAB2221AADB", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CCA211ACA000", 
x"CCAB2111ACAB", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CAB221ACB000", 
x"CCAB2141ACBB", 
x"CAB221ACB000", 
x"CAB221ACB000", 
x"CCA111CCA000", 
x"CCAB2121ACCB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCAB2121ACDB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CCA211ACA000", 
x"B1B000000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCA111CCA000", 
x"CAB121CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CCAB1211CAAB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CCAB1221CACB", 
x"CC11CC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAB1221CADB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CCAB1411CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CA11CA000000", 
x"CCAB1421CBCB", 
x"CC11CC000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CCAB1421CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CCA111CCA000", 
x"CCAB1111CCAB", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CAB121CCB000", 
x"CCAB1141CCBB", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CCA111CCA000", 
x"CCAB1121CCCB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAB1121CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCAB1411CDAB", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CA11CA000000", 
x"CCAB1421CDCB", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAB1421CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB211AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CCA211ACA000", 
x"CAB221ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CAB221ADB000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21DB000000", 
x"CC11CC000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CCA111CCA000", 
x"CAB121CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CAB121CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CCAC2211AAAC", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"CAC211AAC000", 
x"CC11CC000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCAC2111ACAC", 
x"CCA211ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CCAC2141ACBC", 
x"AC11AC000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CCAC2121ACDC", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"AC11AC000000", 
x"CC11CC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAC1211CAAC", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAC1241CABC", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAC1221CADC", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCAC1411CBAC", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAC1441CBBC", 
x"C1C000000000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CC11CC000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAC1421CBDC", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCAC1111CCAC", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAC1141CCBC", 
x"CC11CC000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CCAC1121CCCC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAC1121CCDC", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CCAC1411CDAC", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAC1441CDBC", 
x"C1C000000000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CC11CC000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAC1421CDDC", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"AC11AC000000", 
x"CC11CC000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CCAD2211AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCAD2111ACAD", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAD2141ACBD", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAD2121ACDD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CA11CA000000", 
x"AD11AD000000", 
x"CC11CC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCAD1211CAAD", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CC11CC000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCAD1411CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAD1441CBBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCAD1421CBCD", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCAD1111CCAD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAD1141CCBD", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAD1121CCCD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCAD1121CCDD", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CCAD1411CDAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCAD1441CDBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCAD1421CDCD", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCBA2211AABA", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"BA11BA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CCBA2141ACAA", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCBA2111ACBA", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCBA2141ACDA", 
x"CCB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CCB211ACB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CCB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CCB221AAB000", 
x"CBA141CAA000", 
x"CBA141CAA000", 
x"CCBA1211CABA", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCBA1241CACA", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCBA1241CADA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CCBA1411CBBA", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CCBA1141CCAA", 
x"CCB121CAB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCBA1111CCBA", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCBA1141CCCA", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCBA1141CCDA", 
x"CC3B1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CBA141CDA000", 
x"CB21AB000000", 
x"CBA141CDA000", 
x"CBA141CDA000", 
x"CCBA1411CDBA", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCBA1441CDDA", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"A1A000000000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CBA141CDA000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"A1A000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"CCBB2211AABB", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB3B2141ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB3B2141ABDB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CCBB2111ACBB", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCBB2141ACDB", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"CBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CBB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCBB1241CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCBB1211CABB", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCBB1241CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB3B1141CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB3B1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCBB1141CCAB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCBB1111CCBB", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCBB1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCBB1441CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"CCBB1411CDBB", 
x"CBB141CDB000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCBB1441CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCBC2211AABC", 
x"CCB221AAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB11CB000000", 
x"CBC211ABC000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCBC2141ACAC", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCBC2111ACBC", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCBC2141ACDC", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CCB121CAB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CCB111CCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB221AAB000", 
x"CCBC1241CAAC", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCBC1211CABC", 
x"CCB121CAB000", 
x"CBC141CAC000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCBC1241CADC", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CCBC1411CBBC", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB121CAB000", 
x"CCBC1141CCAC", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCBC1111CCBC", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCBC1141CCCC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC3B1141CCDB", 
x"CCBC1141CCDC", 
x"CC11CC000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CCBC1441CDAC", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCBC1411CDBC", 
x"CCB141CDB000", 
x"CBC141CDC000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CCBC1441CDDC", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCBD2211AABD", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"CCBD2141ACAD", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCBD2111ACBD", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"CCBD2141ACDD", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"B1B000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CCB141CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"CB11CB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"CCBD1241CAAD", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCBD1211CABD", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCBD1241CACD", 
x"CBD141CAD000", 
x"B1B000000000", 
x"CBD141CAD000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CCBD1411CBBD", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CC11CC000000", 
x"CCB121CAB000", 
x"CC11CC000000", 
x"CCBD1141CCAD", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCBD1111CCBD", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CCBD1141CCCD", 
x"CC11CC000000", 
x"CC3B1141CCDB", 
x"CC11CC000000", 
x"CCBD1141CCDD", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCBD1441CDAD", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCBD1411CDBD", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"B1B000000000", 
x"CBD141CDD000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"C1C000000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCCA2211AACA", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCC121CAC000", 
x"CCA211ACA000", 
x"CCCA2141ACBA", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CCCA2111ACCA", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CCCA2141ACDA", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCC121CAC000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCCA1211CACA", 
x"CCC121CAC000", 
x"CC11CC000000", 
x"CCC121CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCA1411CBCA", 
x"CCC141CBC000", 
x"CC11CC000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCCA1141CCBA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCA1111CCCA", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCCA1141CCDA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCA1411CDCA", 
x"CCC141CDC000", 
x"CC11CC000000", 
x"CCC141CDC000", 
x"CCCA1441CDDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"CCA211ACA000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCC121CAC000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"CCCB2221AAAB", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"CCCB2211AACB", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCCB2121ACAB", 
x"CCC121CAC000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"CCCB2111ACCB", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCCB2141ACDB", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"CCC121CAC000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CCB141CDB000", 
x"CCC141CDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCCB1221CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCC121CAC000", 
x"CCCB1211CACB", 
x"CC11CC000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"CCCB1241CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CCCB1411CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCCB1121CCAB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCC111CCC000", 
x"CCCB1111CCCB", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CCCB1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCCB1421CDAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCC141CDC000", 
x"CCCB1411CDCB", 
x"CC11CC000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"CCCB1441CDDB", 
x"C1C000000000", 
x"C1C000000000", 
x"000000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1221CAAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1241CABC", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCC121CAC000", 
x"CCCC1211CACC", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1241CADC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1421CBAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1441CBBC", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCC141CBC000", 
x"CCCC1411CBCC", 
x"CCC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1441CBDC", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCC1121CCAC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCC1141CCBC", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCCC1111CCCC", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCC1141CCDC", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1421CDAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1441CDBC", 
x"C1C000000000", 
x"CCC141CDC000", 
x"CCC141CDC000", 
x"CCCC1411CDCC", 
x"CCC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCC1441CDDC", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCCD2221AAAD", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCCD2211AACD", 
x"CCD221AAD000", 
x"CCD221AAD000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCCD2121ACAD", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCCD2141ACBD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCCD2111ACCD", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CCC141CDC000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCC141CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCD1221CAAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCD1241CABD", 
x"CCC121CAC000", 
x"CCC121CAC000", 
x"CC11CC000000", 
x"CCCD1211CACD", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCCD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCC141CBC000", 
x"CC11CC000000", 
x"CCCD1411CBCD", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCD1121CCAD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCCD1141CCBD", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCCD1111CCCD", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCC141CDC000", 
x"CCC141CDC000", 
x"CC11CC000000", 
x"CCCD1411CDCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCC141CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCDA2211AADA", 
x"CCD221AAD000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CCDA2121ACAA", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"CCDA2141ACBA", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCDA2111ACDA", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CCDA1241CABA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDA1241CACA", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCDA1211CADA", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CCDA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CCDA1411CBDA", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCDA1121CCAA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDA1141CCBA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDA1141CCCA", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCDA1111CCDA", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CCDA1411CDDA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"CCDB2221AAAB", 
x"C1C000000000", 
x"CCD221AAD000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD221AAD000", 
x"CCDB2211AADB", 
x"C1C000000000", 
x"CCD221AAD000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CCDB2121ACAB", 
x"C1C000000000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"CCDB2141ACBB", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCDB1141CC3B", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD211ACD000", 
x"CCDB2111ACDB", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"B1B000000000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCDB1141CC3B", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCDB1221CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"CCDB1241CACB", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD121CAD000", 
x"CCDB1211CADB", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"CCDB1421CBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"CCDB1441CBCB", 
x"CC11CC000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CCDB1411CBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCDB1121CCAB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDB1141CC3B", 
x"CCDB1141CCBB", 
x"CCDB1141CC3B", 
x"CCDB1141CC3B", 
x"CC11CC000000", 
x"CCDB1141CCCB", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCDB1111CCDB", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CCDB1421CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD3B1141CDCB", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCDB1411CDDB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CCDB1141CC3B", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD221AAD000", 
x"CCD221AAD000", 
x"CCDC2211AADC", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC2121ACAC", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC2141ACBC", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CCDC2111ACDC", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"DC11DC000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC1221CAAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC1241CABC", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CC11CC000000", 
x"CDC121CAC000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCDC1211CADC", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC1421CBAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDC1441CBBC", 
x"C1C000000000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CC11CC000000", 
x"CDC141CBC000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"CCDC1411CBDC", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDC1121CCAC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDC1141CCBC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDC1141CCCC", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCDC1111CCDC", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCDC1421CDAC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CCDC1411CDDC", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"CDC211ADC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC121CAC000", 
x"CCD121CAD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CBC000", 
x"DC11DC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD221AAD000", 
x"CCD221AAD000", 
x"C1C000000000", 
x"CCDD2211AADD", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDD2141ACBD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"CCDD2111ACDD", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CCD221AAD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDD1221CAAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDD1241CABD", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"CCDD1211CADD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCDD1441CBBD", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CCDD1411CBDD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDD1121CCAD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCDD1141CCBD", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCDD1111CCDD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAA2111ADAA", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDAA2141ADBA", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDAA2121ADCA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDAA1211CAAA", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDAA1241CABA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAA1221CACA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDAA1221CADA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAA1411CBAA", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDAA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAA1421CBCA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDAA1421CBDA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAA1411CCAA", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAA1111CDAA", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDAA1141CDBA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAA1121CDCA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAA1121CDDA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AA11AA000000", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"CDAB2211AAAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"C1C000000000", 
x"CDAB2221AACB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CDAB2221AADB", 
x"C1C000000000", 
x"CD21AD000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"CDA121CAA000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"CDA141CCA000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDAB1141CD3B", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CDAB2111ADAB", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"DAB221ADB000", 
x"CDAB2141ADBB", 
x"DAB221ADB000", 
x"DAB221ADB000", 
x"C1C000000000", 
x"CDAB2121ADCB", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"CDAB2121ADDB", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDA121CAA000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDAB1141CD3B", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDA121CAA000", 
x"CDAB1211CAAB", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"AB11AB000000", 
x"CDAB1241CABB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"CDAB1221CACB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CDAB1221CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"CDAB1411CBAB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CDAB1441CBBB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CDAB1421CBCB", 
x"AB21CB000000", 
x"CD11CD000000", 
x"AB21CB000000", 
x"CDAB1421CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CDA121CAA000", 
x"CDAB1411CCAB", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"AB21CB000000", 
x"CDAB1441CCBB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CDA141CCA000", 
x"CDAB1421CCCB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDAB1421CCDB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDAB1111CDAB", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDAB1141CD3B", 
x"CDAB1141CDBB", 
x"CDAB1141CD3B", 
x"CDAB1141CD3B", 
x"CD11CD000000", 
x"CDAB1121CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAB1121CDDB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DAB211AAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA3B1141DACB", 
x"DA11DA000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA3B1141DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CD11CD000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CDA121CAA000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"CDA141CCA000", 
x"AB21CB000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDAB1141CD3B", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"C1C000000000", 
x"DAB121DCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"C1C000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CDAC2211AAAC", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDAC2111ADAC", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDAC2141ADBC", 
x"CD21AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAC2121ADCC", 
x"CD11CD000000", 
x"DA11DA000000", 
x"CD21AD000000", 
x"CDAC2121ADDC", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC121DCC000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDAC1211CAAC", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAC1241CABC", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CDAC1221CACC", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"C1C000000000", 
x"CDAC1221CADC", 
x"C1C000000000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDAC1411CBAC", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAC1441CBBC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAC1421CBCC", 
x"CD11CD000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"CDAC1421CBDC", 
x"C1C000000000", 
x"CDA121CAA000", 
x"CDA141CCA000", 
x"CDAC1411CCAC", 
x"CDA141CCA000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"CDAC1441CCBC", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"CDAC1421CCCC", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CDAC1421CCDC", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDAC1111CDAC", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAC1141CDBC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAC1121CDCC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAC1121CDDC", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CDAD2211AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDAD2111ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DAD141DBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DAD121DDD000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDAD1211CAAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAD1241CABD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA211ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"CDAD1221CADD", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDAD1411CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAD1441CBBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAD1421CBDD", 
x"CDA121CAA000", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"CDAD1411CCAD", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDAD1441CCBD", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDAD1111CDAD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAD1141CDBD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAD1121CDCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDAD1121CDDD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CD11CD000000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DAD141DBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"A1A000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDBA2211AABA", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"BA11BA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBA2141ADAA", 
x"DB21AB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDBA2111ADBA", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDBA2141ADDA", 
x"DB11DB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CDB211ADB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDBA1241CAAA", 
x"CDB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDBA1211CABA", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDBA1241CACA", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDBA1241CADA", 
x"CDB211ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"CDBA1411CBBA", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDBA1441CCAA", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDBA1411CCBA", 
x"CDB141CBB000", 
x"CDB141CCB000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBA1141CDAA", 
x"CD3B1141CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBA1111CDBA", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDBA1141CDCA", 
x"CD3B1141CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBA1141CDDA", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DBA141DAA000", 
x"CDB221AAB000", 
x"DBA141DAA000", 
x"DBA141DAA000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DBA141DDA000", 
x"DB21AB000000", 
x"DBA141DDA000", 
x"DBA141DDA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB221AAB000", 
x"CDBB2211AABB", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"DB3B2141ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB3B2141ABCB", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDBB2141ADAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"CDBB2111ADBB", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CDBB2141ADCB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"DBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"CDB141CCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DBB141DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DBB141DCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDBB1241CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDBB1211CABB", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"CDBB1241CACB", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"CDBB1241CADB", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDBB1441CBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"CDBB1411CBBB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDBB1441CBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"CDBB1411CCBB", 
x"CDB141CCB000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBB1141CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDBB1111CDBB", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CDBB1141CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDBB1141CDDB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"DBB211ABB000", 
x"DBB141DAB000", 
x"DBB141DAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB3B1141DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB3B1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB3B1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBB141DCB000", 
x"BB11BB000000", 
x"DBB141DCB000", 
x"DBB141DCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBB141DCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"000000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDBC2211AABC", 
x"CDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"CDBC2141ADAC", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDBC2111ADBC", 
x"CDB211ADB000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDBC2141ADCC", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB11DB000000", 
x"CDBC2141ADDC", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CDB121CAB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CDB111CDB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB221AAB000", 
x"CDBC1241CAAC", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDBC1211CABC", 
x"CDB121CAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDBC1241CACC", 
x"CD11CD000000", 
x"C1C000000000", 
x"CDB211ADB000", 
x"CDBC1241CADC", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDBC1441CBAC", 
x"B1B000000000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDBC1411CBBC", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"CDBC1441CBDC", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDBC1441CCAC", 
x"C1C000000000", 
x"CDB141CCB000", 
x"CDB141CBB000", 
x"CDBC1411CCBC", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"CDBC1441CCCC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD3B1141CDAB", 
x"CDBC1141CDAC", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDBC1111CDBC", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD3B1141CDCB", 
x"CDBC1141CDCC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CDBC1141CDDC", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"CDB141CCB000", 
x"DBC141DCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"B1B000000000", 
x"DBC141DDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"000000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDBD2211AABD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DBD211ABD000", 
x"DB11DB000000", 
x"DBD211ABD000", 
x"DBD211ABD000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDBD2141ADAD", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDBD2111ADBD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CDBD2141ADDD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CDB141CCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"CDBD1241CAAD", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDBD1211CABD", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"CDB211ADB000", 
x"C1C000000000", 
x"CDBD1241CADD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDBD1411CBBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"CDBD1441CCAD", 
x"CDB141CCB000", 
x"CDB141CBB000", 
x"CDB141CCB000", 
x"CDBD1411CCBD", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD3B1141CDAB", 
x"CD11CD000000", 
x"CDBD1141CDAD", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDBD1111CDBD", 
x"CD11CD000000", 
x"CD3B1141CDCB", 
x"CD11CD000000", 
x"CDBD1141CDCD", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CDBD1141CDDD", 
x"D1D000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DBD141DAD000", 
x"CDB211ADB000", 
x"DBD141DAD000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DBD141DDD000", 
x"DB11DB000000", 
x"DBD141DDD000", 
x"DBD141DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CDCA2211AACA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"CDC121CAC000", 
x"DCA211ACA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CDCA2121ADAA", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDCA2141ADBA", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"CDCA2111ADCA", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CD11CD000000", 
x"CDCA2141ADDA", 
x"CD21AD000000", 
x"DC11DC000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CDC121CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CDCA1211CACA", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CDC211ADC000", 
x"CA11CA000000", 
x"CDCA1421CBAA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCA1411CBCA", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDCA1441CBDA", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CDC121CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CDCA1411CCCA", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CDCA1121CDAA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCA1141CDBA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCA1111CDCA", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDCA1141CDDA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"CDC211ADC000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"DCA141DBA000", 
x"C1C000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CBC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"DCA121DAA000", 
x"DCA141DDA000", 
x"C1C000000000", 
x"DCA141DDA000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"CDCB2221AAAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"CDCB2211AACB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CD11CD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCB1141CD3B", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDCB2121ADAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"CDCB2141ADBB", 
x"B1B000000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"CDCB2111ADCB", 
x"CDC211ADC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDCB2141ADDB", 
x"DC11DC000000", 
x"CD21AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDC121CAC000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCB1141CD3B", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDCB1221CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CDCB1241CABB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CDC121CAC000", 
x"CDCB1211CACB", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"CDCB1241CADB", 
x"CDC211ADC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CDCB1411CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CDCB1421CCAB", 
x"CDC121CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CDC141CCC000", 
x"CDCB1411CCCB", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CDCB1141CD3B", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCB1121CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCB1141CD3B", 
x"CDCB1141CDBB", 
x"CDCB1141CD3B", 
x"CDCB1141CD3B", 
x"CDC111CDC000", 
x"CDCB1111CDCB", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CDCB1141CDDB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"CDC211ADC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"CDC121CAC000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCB1141CD3B", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC2211AACC", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDCC2121ADAC", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDCC2141ADBC", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CDCC2111ADCC", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"DC11DC000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC211ACC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC1221CAAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC1241CABC", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDCC1211CACC", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC1241CADC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC1421CBAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCC1441CBBC", 
x"C1C000000000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDCC1411CBCC", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CDC121CAC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CDCC1411CCCC", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CDC111CDC000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCC1121CDAC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCC1141CDBC", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDCC1111CDCC", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCC1141CDDC", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"DCC121DAC000", 
x"DCC211ACC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"CDC211ADC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"DCC141DBC000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC121CAC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CBC000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDCD2121ADAD", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDCD2141ADBD", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CDC211ADC000", 
x"CDCD2111ADCD", 
x"CD21AD000000", 
x"CD21AD000000", 
x"DC11DC000000", 
x"CDCD2141ADDD", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDC211ADC000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCD1221CAAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCD1241CABD", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDCD1211CACD", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC211ADC000", 
x"CDCD1241CADD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDCD1441CBBD", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDCD1411CBCD", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"CDCD1441CBDD", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CDCD1421CCAD", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDCD1411CCCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCD1121CDAD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCD1141CDBD", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDCD1111CDCD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDCD1141CDDD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCD121DAD000", 
x"DCD121DAD000", 
x"CDC211ADC000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCD141DBD000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC121CAC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CBC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"CDC111CDC000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD141DDD000", 
x"DCD141DDD000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDDA2211AADA", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"CDDA2141ADBA", 
x"CD21AD000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDDA2111ADDA", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DDA211ADA000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CDDA1221CAAA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDA1241CABA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDA1241CACA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDDA1211CADA", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDDA1421CBAA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDA1441CBBA", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDA1441CBCA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDDA1411CBDA", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDDA1421CCAA", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"CDDA1441CCBA", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"CDDA1441CCCA", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDDA1411CCDA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDDA1121CDAA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDA1141CDBA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDA1141CDCA", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDA1111CDDA", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"CDD211ADD000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CD11CD000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"CDDB2221AAAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CDDB2211AADB", 
x"C1C000000000", 
x"CDD211ADD000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD21AD000000", 
x"CDDB2121ADAB", 
x"C1C000000000", 
x"CD21AD000000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"C1C000000000", 
x"CDDB2141ADCB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD211ADD000", 
x"CDDB2111ADDB", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDDB1221CAAB", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"CDDB1241CABB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDDB1241CACB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD121CAD000", 
x"CDDB1211CADB", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"CDDB1421CBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDDB1441CBBB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDDB1441CBCB", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CDDB1411CBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDDB1421CCAB", 
x"C1C000000000", 
x"CDD121CAD000", 
x"B1B000000000", 
x"CDDB1441CCBB", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDDB1441CCCB", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDB1411CCDB", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD11CD000000", 
x"CDDB1121CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CDDB1141CDBB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CDDB1141CDCB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDDB1111CDDB", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DD11DD000000", 
x"DDB121DAB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDB141DCB000", 
x"DD11DD000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDDC2211AADC", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDDC2121ADAC", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"CDDC2141ADBC", 
x"CD21AD000000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"CD11CD000000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDDC2111ADDC", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"DDC211ADC000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1221CAAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1241CABC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1241CACC", 
x"CD11CD000000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDDC1211CADC", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1421CBAC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1441CBBC", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1441CBCC", 
x"CD11CD000000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDDC1411CBDC", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1421CCAC", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1441CCBC", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDC1441CCCC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDC1411CCDC", 
x"CDD111CDD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDC1121CDAC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDC1141CDBC", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDC1141CDCC", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDDC1111CDDC", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"CDD211ADD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CDD121CAD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC121DAC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC141DBC000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDDD2121ADAD", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDDD2141ADBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"CDDD2111ADDD", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD21AD000000", 
x"CD21AD000000", 
x"C1C000000000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"CD21AD000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DDD141DBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDD1221CAAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDD1241CABD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"CDDD1211CADD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDD1421CBAD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDDD1441CBBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"CDDD1411CBDD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDD1121CDAD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDD1141CDBD", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDDD1141CDCD", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDDD1111CDDD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"CDD211ADD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDD111CDD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"CD11CD000000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DA11DA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AAA111AAA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AAA121ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAA1111DAAA", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAAA1141DABA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAA1121DACA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAA1121DADA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAA1411DBAA", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"DAAA1441DBBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAA1421DBCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAA1211DCAA", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAAA1241DCBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAA1221DCCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"DAAB2111AAAB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"DAAB2121AACB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DA11DA000000", 
x"DAAB2121AADB", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AA11AA000000", 
x"DAAB2211ACAB", 
x"A1A000000000", 
x"D1D000000000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"DAAB2221ACCB", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAAB2221ACDB", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DAAB2211ADAB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"AAB121ADB000", 
x"DAA121DCA000", 
x"DAAB2221ADCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAAB2221ADDB", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"AAB111AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"AAB121ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB121ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AAB211CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAA111DAA000", 
x"AAB211DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AAB111AAB000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"AAB121ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AAB121ADB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AA11AA000000", 
x"AAB211CAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"AAB221CCB000", 
x"A1A000000000", 
x"AAB221CCB000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AAB221CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"AAB211DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"AAB221CDB000", 
x"DAA121DCA000", 
x"AAB221DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AAB221DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DAAB1111DAAB", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"AAB211DAB000", 
x"DAAB1141DABB", 
x"AAB211DAB000", 
x"AAB211DAB000", 
x"DA11DA000000", 
x"DAAB1121DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAB1121DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DAAB1411DBAB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAAB1441DBBB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAAB1421DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAAB1421DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAA121DCA000", 
x"DAAB1211DCAB", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"AAB221DCB000", 
x"DAAB1241DCBB", 
x"AAB221DCB000", 
x"AAB221DCB000", 
x"D1D000000000", 
x"DAAB1221DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAAB1221DCDB", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DAAB1211DDAB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AAB221DDB000", 
x"DAAB1241DDBB", 
x"AAB221DDB000", 
x"AAB221DDB000", 
x"DAA121DCA000", 
x"DAAB1221DDCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAAB1221DDDB", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DAAC2111AAAC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DAAC2141AABC", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"AAC111AAC000", 
x"DA11DA000000", 
x"AA11AA000000", 
x"DAAC2121AADC", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"AAC141ABC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DAAC2211ADAC", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"AAC121ADC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAAC2221ADDC", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAC141ABC000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AAC121ADC000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"AAC211DAC000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AAC221DDC000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAC111AAC000", 
x"AA11AA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AAC141ABC000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"AAC211CAC000", 
x"DA11DA000000", 
x"C1C000000000", 
x"AAC121ADC000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AA11AA000000", 
x"C1C000000000", 
x"AAC211CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"AAC211DAC000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAA121DCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAAC1111DAAC", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAC1141DABC", 
x"DA11DA000000", 
x"AAC211DAC000", 
x"AAC211DAC000", 
x"DAAC1121DACC", 
x"AAC211DAC000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAC1121DADC", 
x"DA11DA000000", 
x"AA11AA000000", 
x"DAA141DBA000", 
x"DAAC1411DBAC", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAC1441DBBC", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAAC1421DBCC", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAAC1421DBDC", 
x"D1D000000000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAAC1211DCAC", 
x"DAA121DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAAC1241DCBC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAAC1221DCCC", 
x"AC21DC000000", 
x"DA11DA000000", 
x"AC21DC000000", 
x"DAAC1221DCDC", 
x"AC21DC000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DAAC1211DDAC", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"DAAC1241DDBC", 
x"D1D000000000", 
x"DAA121DCA000", 
x"AAC221DDC000", 
x"DAAC1221DDCC", 
x"AAC221DDC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAAC1221DDDC", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DAAD2111AAAD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AAD111AAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AAD141ABD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAAD2211ACAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"AAD121ACD000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DAA121DCA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AAD111AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD121ACD000", 
x"DA11DA000000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AAD211CAD000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AAD211CAD000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAAD1111DAAD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAD1141DABD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAD1121DACD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAD1121DADD", 
x"AA11AA000000", 
x"DAA141DBA000", 
x"DAA141DBA000", 
x"DAAD1411DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1441DBBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1421DBCD", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1421DBDD", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAAD1211DCAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1241DCBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1221DCCD", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1221DCDD", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAAD1211DDAD", 
x"DAA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1241DDBD", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1221DDCD", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAAD1221DDDD", 
x"ABA141AAA000", 
x"DAB211AAB000", 
x"ABA141AAA000", 
x"ABA141AAA000", 
x"DABA2111AABA", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DABA2141AACA", 
x"DAB221ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"D1D000000000", 
x"D1D000000000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"ABA141ACA000", 
x"DABA2211ACBA", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DABA2211ADBA", 
x"DAB141DBB000", 
x"DAB221ADB000", 
x"DAB221ADB000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"DAB211AAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"AB11AB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA211CBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA211DBA000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABA141AAA000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"ABA111ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABA141ACA000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"D1D000000000", 
x"D1D000000000", 
x"ABA211CBA000", 
x"AB11AB000000", 
x"ABA211CBA000", 
x"ABA211CBA000", 
x"BA11BA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ABA211CBA000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ABA211DBA000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DABA1141DAAA", 
x"DAB211AAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DABA1111DABA", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DABA1141DACA", 
x"DA3B1141DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DABA1141DADA", 
x"DA3B1141DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ABA211DBA000", 
x"AB11AB000000", 
x"ABA211DBA000", 
x"ABA211DBA000", 
x"DABA1411DBBA", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DABA1241DCAA", 
x"AB11AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DABA1211DCBA", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DABA1241DCCA", 
x"AB21CB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DABA1211DDBA", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DABA1241DDCA", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DAB211AAB000", 
x"DABB2111AABB", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"DABB2141AACB", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DABB2141AADB", 
x"D1D000000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"AB3B1141ABAB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB3B1141ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB3B1141ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ABB141ACB000", 
x"DABB2211ACBB", 
x"ABB141ACB000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"ABB141ADB000", 
x"DABB2211ADBB", 
x"ABB141ADB000", 
x"ABB141ADB000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"ABB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"ABB211CBB000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"ABB211DBB000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"ABB111ABB000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"ABB141ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"ABB141ADB000", 
x"D1D000000000", 
x"D1D000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB3B2141CBCB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB3B2141CBDB", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB21CB000000", 
x"ABB211CBB000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DABB1141DAAB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DABB1111DABB", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DABB1141DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DABB1141DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABB211DBB000", 
x"DABB1411DBBB", 
x"ABB211DBB000", 
x"ABB211DBB000", 
x"AB21DB000000", 
x"AB3B2141DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB3B2141DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"DABB1211DCBB", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"DABB1241DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DABB1241DCDB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DABB1211DDBB", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"DABC2141AAAC", 
x"D1D000000000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DABC2111AABC", 
x"DAB211AAB000", 
x"ABC141AAC000", 
x"DAB221ACB000", 
x"ABC141AAC000", 
x"ABC141AAC000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"DABC2141AADC", 
x"D1D000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"BC11BC000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DABC2211ACBC", 
x"DAB221ACB000", 
x"ABC141ACC000", 
x"AB21CB000000", 
x"ABC141ACC000", 
x"ABC141ACC000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"DAB141DBB000", 
x"DABC2211ADBC", 
x"DAB221ADB000", 
x"ABC141ADC000", 
x"DAB121DCB000", 
x"ABC141ADC000", 
x"ABC141ADC000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"ABC211DBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DAB211AAB000", 
x"ABC141AAC000", 
x"C1C000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABC111ABC000", 
x"AB11AB000000", 
x"C1C000000000", 
x"DAB221ACB000", 
x"ABC141ACC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"ABC141ADC000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BC11BC000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABC211CBC000", 
x"AB21CB000000", 
x"C1C000000000", 
x"AB21CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"C1C000000000", 
x"DAB121DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB211AAB000", 
x"DABC1141DAAC", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DABC1111DABC", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA3B1141DACB", 
x"DABC1141DACC", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA3B1141DADB", 
x"DABC1141DADC", 
x"DA11DA000000", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DABC1411DBBC", 
x"DAB141DBB000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"ABC211DBC000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"C1C000000000", 
x"AB11AB000000", 
x"DABC1241DCAC", 
x"C1C000000000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DABC1211DCBC", 
x"DAB121DCB000", 
x"C1C000000000", 
x"AB21CB000000", 
x"DABC1241DCCC", 
x"C1C000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DABC1241DCDC", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DABC1241DDAC", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DABC1211DDBC", 
x"DAB121DDB000", 
x"C1C000000000", 
x"DAB121DCB000", 
x"DABC1241DDCC", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DABC1241DDDC", 
x"D1D000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"DABD2141AAAD", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DABD2111AABD", 
x"A1A000000000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"DABD2141AACD", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"ABD141AAD000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DABD2211ACBD", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"ABD141ACD000", 
x"ABD141ACD000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"DAB141DBB000", 
x"DAB221ADB000", 
x"DABD2211ADBD", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"ABD141ADD000", 
x"ABD141ADD000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ABD211CBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DAB111DAB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DAB121DCB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DAB121DDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"ABD141AAD000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"ABD111ABD000", 
x"A1A000000000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"ABD141ACD000", 
x"DA11DA000000", 
x"DAB221ADB000", 
x"D1D000000000", 
x"ABD141ADD000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"BD11BD000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"ABD211CBD000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DAB211AAB000", 
x"DA11DA000000", 
x"DABD1141DAAD", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DABD1111DABD", 
x"DA11DA000000", 
x"DA3B1141DACB", 
x"DA11DA000000", 
x"DABD1141DACD", 
x"DA11DA000000", 
x"DA3B1141DADB", 
x"DA11DA000000", 
x"DABD1141DADD", 
x"AB21DB000000", 
x"AB11AB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DABD1411DBBD", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"ABD211DBD000", 
x"D1D000000000", 
x"AB11AB000000", 
x"D1D000000000", 
x"DABD1241DCAD", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DABD1211DCBD", 
x"D1D000000000", 
x"AB21CB000000", 
x"D1D000000000", 
x"DABD1241DCCD", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DABD1241DCDD", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DABD1211DDBD", 
x"D1D000000000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"DABD1241DDCD", 
x"DA11DA000000", 
x"DAB121DDB000", 
x"D1D000000000", 
x"DABD1241DDDD", 
x"ACA121AAA000", 
x"ACA121AAA000", 
x"DAC211AAC000", 
x"ACA121AAA000", 
x"DACA2141AABA", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DACA2111AACA", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC221ADC000", 
x"D1D000000000", 
x"ACA141ABA000", 
x"ACA141ABA000", 
x"AC11AC000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DACA2211ADCA", 
x"DAC221ADC000", 
x"DAC121DCC000", 
x"DAC221ADC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"ACA121AAA000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"D1D000000000", 
x"ACA141ABA000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC221ADC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DAC211AAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"ACA111ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"ACA211CCA000", 
x"AC11AC000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACA211CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC141DBC000", 
x"C1C000000000", 
x"ACA211DCA000", 
x"C1C000000000", 
x"DAC121DCC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"DAC121DDC000", 
x"C1C000000000", 
x"DACA1121DAAA", 
x"DA11DA000000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"DACA1141DABA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACA1111DACA", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DACA1141DADA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACA1421DBAA", 
x"D1D000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DACA1441DBBA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DACA1411DBCA", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"ACA211DCA000", 
x"ACA211DCA000", 
x"AC11AC000000", 
x"ACA211DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DACA1211DCCA", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DA11DA000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DACA1241DDBA", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DACA1211DDCA", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"DACB2121AAAB", 
x"DAC211AAC000", 
x"D1D000000000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"ACB121AAB000", 
x"DAC211AAC000", 
x"DACB2111AACB", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"DACB2141AADB", 
x"DAC221ADC000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"CB21AB000000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"ACB141ABB000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"AC11AC000000", 
x"AC3B1141ACAB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"DACB2211ACCB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC3B1141ACDB", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"DACB1141DA3B", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"ACB141ADB000", 
x"DAC221ADC000", 
x"DACB2211ADCB", 
x"DAC121DCC000", 
x"DAC221ADC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"B1B000000000", 
x"ACB121AAB000", 
x"DAC211AAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"ACB141ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"ACB211CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DACB1141DA3B", 
x"DAC111DAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ACB211DCB000", 
x"DAC121DCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB121AAB000", 
x"DAC211AAC000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"ACB141ABB000", 
x"ACB221CAB000", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"ACB111ACB000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"ACB141ADB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"ACB221CAB000", 
x"AC11AC000000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"ACB211CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DACB1141DA3B", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"ACB211DCB000", 
x"DAC121DCC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DACB1121DAAB", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"DACB1141DA3B", 
x"DACB1141DABB", 
x"DACB1141DA3B", 
x"DACB1141DA3B", 
x"DAC111DAC000", 
x"DACB1111DACB", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DACB1141DADB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DACB1421DBAB", 
x"AC11AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DACB1441DBBB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DACB1411DBCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DACB1441DBDB", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"DACB1221DCAB", 
x"AC11AC000000", 
x"AC21DC000000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"ACB211DCB000", 
x"DAC121DCC000", 
x"DACB1211DCCB", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DA11DA000000", 
x"DACB1241DCDB", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"DACB1221DDAB", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DACB1241DDBB", 
x"B1B000000000", 
x"B1B000000000", 
x"DAC121DDC000", 
x"DACB1211DDCB", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DA11DA000000", 
x"DACB1241DDDB", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DACC2141AABC", 
x"D1D000000000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DACC2111AACC", 
x"DAC211AAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DACC2141AADC", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ACC141ABC000", 
x"ACC141ABC000", 
x"CC11CC000000", 
x"ACC141ABC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"ACC141ADC000", 
x"ACC141ADC000", 
x"DACC2211ADCC", 
x"ACC141ADC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ACC141ABC000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"ACC141ADC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"AC21DC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC211AAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACC141ABC000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACC111ACC000", 
x"AC11AC000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"ACC141ADC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC141DBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACC211DCC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"DAC121DDC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACC1121DAAC", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACC1141DABC", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DACC1111DACC", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACC1141DADC", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DACC1441DBBC", 
x"D1D000000000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DACC1411DBCC", 
x"DAC141DBC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DACC1441DBDC", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC11AC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DACC1241DCBC", 
x"AC21DC000000", 
x"ACC211DCC000", 
x"ACC211DCC000", 
x"DACC1211DCCC", 
x"ACC211DCC000", 
x"DA11DA000000", 
x"AC21DC000000", 
x"DACC1241DCDC", 
x"AC21DC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DACC1211DDCC", 
x"DAC121DDC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"DACD2121AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"DACD2141AABD", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DACD2111AACD", 
x"DA11DA000000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"ACD141ABD000", 
x"AC21DC000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"ACD111ACD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DAC221ADC000", 
x"DAC221ADC000", 
x"DAC121DCC000", 
x"DACD2211ADCD", 
x"DA11DA000000", 
x"ACD141ADD000", 
x"DAC121DDC000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"ACD121AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"ACD141ABD000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC221ADC000", 
x"ACD141ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"ACD211DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC211AAC000", 
x"ACD121AAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"ACD111ACD000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"ACD211CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAC111DAC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAC121DCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DAC121DDC000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC211AAC000", 
x"DACD1121DAAD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACD1141DABD", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DACD1111DACD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DACD1141DADD", 
x"D1D000000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"DACD1421DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DACD1441DBBD", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DACD1411DBCD", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"DACD1441DBDD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC11AC000000", 
x"DACD1221DCAD", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DACD1211DCCD", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"ACD211DCD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"DACD1241DDBD", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DACD1211DDCD", 
x"DA11DA000000", 
x"D1D000000000", 
x"DAC121DDC000", 
x"DACD1241DDDD", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"ADA121AAA000", 
x"DAD211AAD000", 
x"DADA2141AABA", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DADA2141AACA", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DADA2111AADA", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"ADA141ABA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"ADA141ACA000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"ADA111ADA000", 
x"DAD111DAD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADA121AAA000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DDD000", 
x"ADA121AAA000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"ADA141ABA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADA141ACA000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"ADA111ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DDD000", 
x"DADA1121DAAA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADA1141DABA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADA1141DACA", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADA1111DADA", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DADA1421DBAA", 
x"D1D000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DADA1441DBBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADA1441DBCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADA1411DBDA", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DADA1221DCAA", 
x"D1D000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DADA1241DCBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADA1241DCCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADA1211DCDA", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DADA1241DDBA", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"DADA1241DDCA", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DADA1211DDDA", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"A1A000000000", 
x"DADB2121AAAB", 
x"A1A000000000", 
x"DAD211AAD000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"DADB2141AACB", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DADB2111AADB", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"ADB141ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"DADB2221ACAB", 
x"A1A000000000", 
x"AD11AD000000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DADB2211ACDB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DADB1141DA3B", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD3B1141ADCB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DA11DA000000", 
x"DADB2211ADDB", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"ADB121AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ABB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB141ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB111ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211CDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DADB1141DA3B", 
x"B1B000000000", 
x"DAD111DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"ADB211DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB121AAB000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"ADB221CAB000", 
x"ADB141ABB000", 
x"ADB221CAB000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"ADB141ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"ADB111ADB000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"ADB221CAB000", 
x"A1A000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"ADB211CDB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DADB1141DA3B", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"ADB211CDB000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"ADB211DDB000", 
x"D1D000000000", 
x"DAD121DDD000", 
x"DA11DA000000", 
x"DADB1121DAAB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADB1141DA3B", 
x"DADB1141DABB", 
x"DADB1141DA3B", 
x"DADB1141DA3B", 
x"DA11DA000000", 
x"DADB1141DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DADB1111DADB", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DADB1411DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DADB1221DCAB", 
x"D1D000000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"DADB1241DCBB", 
x"B1B000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DADB1241DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DADB1211DCDB", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"DADB1221DDAB", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"ADB211DDB000", 
x"D1D000000000", 
x"DADB1241DDCB", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"DADB1211DDDB", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DADC2121AAAC", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DADC2141AABC", 
x"D1D000000000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"ADC121AAC000", 
x"DA11DA000000", 
x"DAD211AAD000", 
x"DADC2111AADC", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"ADC141ABC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"ADC141ACC000", 
x"DA11DA000000", 
x"DC21AC000000", 
x"DADC2211ACDC", 
x"DC21AC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"ADC111ADC000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"DADC2211ADDC", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC121AAC000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADC141ABC000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"ADC141ACC000", 
x"DC21AC000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DAD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"ADC211DDC000", 
x"DAD121DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC121AAC000", 
x"DAD211AAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC141ABC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"ADC141ACC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"ADC111ADC000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"ADC211CDC000", 
x"C1C000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAD141DBD000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"ADC211CDC000", 
x"DA11DA000000", 
x"C1C000000000", 
x"ADC211DDC000", 
x"DAD121DDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADC1121DAAC", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADC1141DABC", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADC1141DACC", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DADC1111DADC", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADC1421DBAC", 
x"AD11AD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADC1441DBBC", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DADC1441DBCC", 
x"C1C000000000", 
x"DA11DA000000", 
x"DAD141DBD000", 
x"DADC1411DBDC", 
x"DAD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DADC1211DCDC", 
x"DC11DC000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADC1221DDAC", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADC1241DDBC", 
x"DAD141DBD000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"ADC211DDC000", 
x"DA11DA000000", 
x"DAD121DDD000", 
x"DADC1211DDDC", 
x"DAD121DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DADD2141AABD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DADD2141AACD", 
x"DA11DA000000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"DADD2111AADD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"ADD141ABD000", 
x"ADD141ABD000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"ADD141ACD000", 
x"ADD141ACD000", 
x"DADD2211ACDD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADD211CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DAD121DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ABD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"ADD141ACD000", 
x"DA11DA000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"ADD111ADD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"ADD211CDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"ADD211CDD000", 
x"ADD211CDD000", 
x"DAD121DDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADD1121DAAD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADD1141DABD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DADD1141DACD", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DADD1111DADD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADD1441DBBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADD1441DBCD", 
x"DA11DA000000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DADD1411DBDD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADD1241DCBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DADD1241DCCD", 
x"DA11DA000000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DADD1211DCDD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DAD121DCD000", 
x"DA11DA000000", 
x"DAD121DDD000", 
x"DAD121DDD000", 
x"DADD1211DDDD", 
x"AA11AA000000", 
x"DB21AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AA11AA000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DB11DB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DBAA2111ABAA", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"BA11BA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAA2121ABCA", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAA2121ABDA", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AA11AA000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DB11DB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BAA121BCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"BAA121BDA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"DB21AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BAA111BAA000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAA121BDA000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AA11AA000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBAA1411DAAA", 
x"DB21AB000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAA1421DACA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBAA1421DADA", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBAA1111DBAA", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBAA1141DBBA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAA1121DBCA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAA1121DBDA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAA1411DCAA", 
x"DB21AB000000", 
x"DBA141DCA000", 
x"DBA141DCA000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBAA1421DCCA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBAA1421DCDA", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBAA1411DDAA", 
x"DB21AB000000", 
x"DBA141DDA000", 
x"DBA141DDA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAA1421DDCA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"DBAB2111ABAB", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"BA11BA000000", 
x"DBAB2141ABBB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"DBAB2121ABCB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"DBAB2121ABDB", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"AB11AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DBAB1141DB3B", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B3AB1411BAAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA3B1141BACB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA3B1141BADB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB121BCB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"BAB121BDB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B3AB1411BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B3AB1421BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AB1411BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B3AB1421BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BAB111BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAB141BBB000", 
x"BAB141B3B000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"BAB121BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAB121BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"AB11AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DBAB1141DB3B", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"DBAB1411DAAB", 
x"DBA141DAA000", 
x"DBA141DAA000", 
x"DBA211ABA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"D1D000000000", 
x"DBAB1421DACB", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DBAB1111DBAB", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBAB1141DB3B", 
x"DBAB1141DBBB", 
x"DBAB1141DB3B", 
x"DBAB1141DB3B", 
x"DB11DB000000", 
x"DBAB1121DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAB1121DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"DBAB1411DCAB", 
x"DBA141DCA000", 
x"DBA141DCA000", 
x"BA11BA000000", 
x"BAB141B3B000", 
x"B1B000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBAB1421DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DBAB1411DDAB", 
x"DBA141DDA000", 
x"DBA141DDA000", 
x"DBA111DBA000", 
x"DBAB1141DB3B", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"DBAB1421DDCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBAC2111ABAC", 
x"DBA211ABA000", 
x"BA11BA000000", 
x"DB21AB000000", 
x"DBAC2141ABBC", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAC2121ABCC", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DBAC2121ABDC", 
x"DB21AB000000", 
x"AC11AC000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DB11DB000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DBA141DAA000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"DB11DB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"BAC141BBC000", 
x"BAC121BCC000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BCAC", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AC1411BDAC", 
x"B1B000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAC111BAC000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"BAC141BBC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAC121BCC000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"BAC121BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBA141DAA000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBA141DAA000", 
x"DB21AB000000", 
x"DBAC1411DAAC", 
x"DBA141DAA000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"AC11AC000000", 
x"B1B000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBAC1421DADC", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBAC1111DBAC", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAC1141DBBC", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAC1121DBCC", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAC1121DBDC", 
x"DB11DB000000", 
x"AC21DC000000", 
x"DB21AB000000", 
x"DBAC1411DCAC", 
x"AC21DC000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"DBAC1421DCCC", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DB11DB000000", 
x"DBAC1421DCDC", 
x"AC21DC000000", 
x"DBA141DDA000", 
x"DB21AB000000", 
x"DBAC1411DDAC", 
x"DBA141DDA000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AC21DC000000", 
x"B1B000000000", 
x"DBAC1421DDCC", 
x"AC21DC000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"DBAC1421DDDC", 
x"D1D000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBAD2111ABAD", 
x"BA11BA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAD2141ABBD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBAD2121ABCD", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DBAD2121ABDD", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DB21AB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"AD11AD000000", 
x"B1B000000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"BAD141BBD000", 
x"DB11DB000000", 
x"BAD141BBD000", 
x"BAD121BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AD1411BCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"DB11DB000000", 
x"BAD121BCD000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3AD1411BDAD", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"DB11DB000000", 
x"BAD121BDD000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DB11DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BAD111BAD000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD141BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BAD121BCD000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"BAD121BDD000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"DB21AB000000", 
x"D1D000000000", 
x"AD11AD000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA141DAA000", 
x"DB21AB000000", 
x"DBA141DAA000", 
x"DBAD1411DAAD", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBAD1421DACD", 
x"AD11AD000000", 
x"DB11DB000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBAD1111DBAD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAD1141DBBD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAD1121DBCD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBAD1121DBDD", 
x"DBA141DCA000", 
x"DB21AB000000", 
x"DBA141DCA000", 
x"DBAD1411DCAD", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBAD1421DCCD", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBAD1421DCDD", 
x"DBA141DDA000", 
x"DB21AB000000", 
x"DBA141DDA000", 
x"DBAD1411DDAD", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBAD1421DDCD", 
x"DBA141DDA000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBAD1421DDDD", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"DB3B2141ABAB", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DBBA2111ABBA", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBBA2141ABCA", 
x"DB3B2141ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBBA2141ABDA", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B3BA1411BABA", 
x"DBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DB11DB000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"BBA141BCA000", 
x"B3BA1411BCBA", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"DBB141DAB000", 
x"BBA141BDA000", 
x"BBA141BDA000", 
x"B3BA1411BDBA", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DBB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B3B141BAB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BBA111BBA000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBA141BCA000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBA141BDA000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1441DAAA", 
x"DB21AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1411DABA", 
x"DBB211ABB000", 
x"DBB141DAB000", 
x"DBB141DAB000", 
x"DBBA1441DACA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1441DADA", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1141DBAA", 
x"DB3B1141DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBBA1111DBBA", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBBA1141DBCA", 
x"DB3B1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBBA1141DBDA", 
x"DB3B1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBBA1441DCAA", 
x"DB21AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1411DCBA", 
x"BB11BB000000", 
x"DBB141DCB000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1441DCDA", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1441DDAA", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1411DDBA", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBBA1441DDCA", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBA1441DDDA", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBBB2141ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DBBB2111ABBB", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DBBB2141ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBBB2141ABDB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3BB1441BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B3BB1411BABB", 
x"BBB141BAB000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"BB3B1441BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB3B1141BBAB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB3B1141BBCB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB3B1141BBDB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B3BB1441BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B3BB1411BCBB", 
x"BBB141BCB000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B3BB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBB141DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"DBB111DBB000", 
x"BBB141BDB000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"BB3B1441BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BBB141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BBB111BBB000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BBB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBB141BDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBBB1441DAAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"DBBB1411DABB", 
x"DBB141DAB000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"DBBB1441DACB", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBBB1141DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBBB1111DBBB", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DBBB1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBBB1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBBB1441DCAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"DBBB1411DCBB", 
x"DBB141DCB000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB3B2141ABAB", 
x"DBBC2141ABAC", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBBC2111ABBC", 
x"DBB211ABB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DBBC2141ABDC", 
x"DB21AB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBB141DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"DBB211ABB000", 
x"B3BC1411BABC", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BB11BB000000", 
x"B3BC1411BCBC", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DBB141DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"B3BC1411BDBC", 
x"DB11DB000000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"BBC141BAC000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBC111BBC000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"BBC141BDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBB141DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBB141DCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBBC1441DAAC", 
x"D1D000000000", 
x"DBB141DAB000", 
x"DBB211ABB000", 
x"DBBC1411DABC", 
x"DBB141DAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"DBBC1441DACC", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBBC1441DADC", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB3B1141DBAB", 
x"DBBC1141DBAC", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBBC1111DBBC", 
x"DBB111DBB000", 
x"BC11BC000000", 
x"DB3B1141DBCB", 
x"DBBC1141DBCC", 
x"BC11BC000000", 
x"DB11DB000000", 
x"DB3B1141DBDB", 
x"DBBC1141DBDC", 
x"DB11DB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBBC1441DCAC", 
x"C1C000000000", 
x"DBB141DCB000", 
x"BB11BB000000", 
x"DBBC1411DCBC", 
x"DBB141DCB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBBC1441DCDC", 
x"C1C000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"DBBC1441DDAC", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBBC1411DDBC", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBB141DCB000", 
x"DBBC1441DDCC", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBBC1441DDDC", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB3B2141ABAB", 
x"DB21AB000000", 
x"DBBD2141ABAD", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBBD2111ABBD", 
x"DB21AB000000", 
x"DB3B2141ABCB", 
x"DB21AB000000", 
x"DBBD2141ABCD", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"DBB211ABB000", 
x"B3B141BAB000", 
x"B3BD1411BABD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"DB11DB000000", 
x"BBD141BAD000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3BD1411BCBD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"DB11DB000000", 
x"BBD141BCD000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"B3BD1411BDBD", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"BBD141BAD000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BBD111BBD000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"BBD141BCD000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBBD1441DAAD", 
x"DBB141DAB000", 
x"DBB211ABB000", 
x"DBB141DAB000", 
x"DBBD1411DABD", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBBD1441DACD", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBBD1441DADD", 
x"DB11DB000000", 
x"DB3B1141DBAB", 
x"DB11DB000000", 
x"DBBD1141DBAD", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBBD1111DBBD", 
x"DB11DB000000", 
x"DB3B1141DBCB", 
x"DB11DB000000", 
x"DBBD1141DBCD", 
x"DB11DB000000", 
x"DB3B1141DBDB", 
x"DB11DB000000", 
x"DBBD1141DBDD", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBBD1441DCAD", 
x"DBB141DCB000", 
x"BB11BB000000", 
x"DBB141DCB000", 
x"DBBD1411DCBD", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBBD1441DCDD", 
x"D1D000000000", 
x"DBB141DAB000", 
x"D1D000000000", 
x"DBBD1441DDAD", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DBBD1411DDBD", 
x"D1D000000000", 
x"DBB141DCB000", 
x"D1D000000000", 
x"DBBD1441DDCD", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBBD1441DDDD", 
x"A1A000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBCA2121ABAA", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBCA2141ABBA", 
x"DB21AB000000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"DBCA2111ABCA", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBCA2141ABDA", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"B3CA1411BACA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA121BAA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"BCA141BDA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"B3CA1411BDCA", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"BCA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCA141BBA000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BCA111BCA000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCA141BDA000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"C1C000000000", 
x"DBCA1421DAAA", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBCA1411DACA", 
x"B1B000000000", 
x"DBC141DAC000", 
x"DBC141DAC000", 
x"DBCA1441DADA", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBCA1121DBAA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCA1141DBBA", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DB11DB000000", 
x"DBCA1111DBCA", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBCA1141DBDA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"CA11CA000000", 
x"DB21AB000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DBCA1411DCCA", 
x"B1B000000000", 
x"DBC141DCC000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DBCA1421DDAA", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBCA1411DDCA", 
x"B1B000000000", 
x"DBC141DDC000", 
x"DBC141DDC000", 
x"DBCA1441DDDA", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBCB2141AB3B", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBCB2121ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBCB2141AB3B", 
x"DBCB2141ABBB", 
x"BC11BC000000", 
x"DBCB2141AB3B", 
x"DBC211ABC000", 
x"DBCB2111ABCB", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBCB2141ABDB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBCB1141DB3B", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3CB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"BCB121BAB000", 
x"B1B000000000", 
x"B3CB1411BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141B3B000", 
x"BCB121BAB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB141B3B000", 
x"BCB141BDB000", 
x"BCB141B3B000", 
x"BCB141B3B000", 
x"BC11BC000000", 
x"BC3B1141BCAB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"B3CB1411BCCB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC3B1141BCDB", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B3CB1421BDAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BCB141BDB000", 
x"BCB141BDB000", 
x"DBC111DBC000", 
x"BCB141BDB000", 
x"B1B000000000", 
x"B3CB1411BDCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBCB2141AB3B", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"BCB121BAB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BCB141BBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BCB111BCB000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BCB141BDB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBCB1141DB3B", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBCB1421DAAB", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBCB2141AB3B", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"DBCB1411DACB", 
x"DBC141DAC000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBCB1121DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCB1141DB3B", 
x"DBCB1141DBBB", 
x"DBCB1141DB3B", 
x"DBCB1141DB3B", 
x"DBC111DBC000", 
x"DBCB1111DBCB", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBCB1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBCB1421DCAB", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"DBC141DCC000", 
x"DBCB1411DCCB", 
x"DBC141DCC000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DBCB1421DDAB", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBCB1141DB3B", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"DBCB1411DDCB", 
x"DBC141DDC000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBCC2121ABAC", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBCC2111ABCC", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DBCC2141ABDC", 
x"DB21AB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"BCC141BDC000", 
x"BCC141BDC000", 
x"B3CC1411BDCC", 
x"BCC141BDC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCC111BCC000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"BCC141BDC000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"BC11BC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"DB11DB000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBCC1421DAAC", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"B1B000000000", 
x"DBCC1411DACC", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBCC1441DADC", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCC1121DBAC", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCC1141DBBC", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBCC1111DBCC", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCC1141DBDC", 
x"DB11DB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DBCC1421DCAC", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"DBCC1411DCCC", 
x"CC11CC000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"B1B000000000", 
x"DBCC1411DDCC", 
x"DBC141DDC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"000000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBCD2121ABAD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BC11BC000000", 
x"DBCD2141ABBD", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBCD2111ABCD", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DBCD2141ABDD", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BACD", 
x"BCD121BAD000", 
x"DB11DB000000", 
x"BCD121BAD000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD141BBD000", 
x"DB11DB000000", 
x"BCD141BBD000", 
x"BCD141BDD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3CD1411BDCD", 
x"BCD141BDD000", 
x"DB11DB000000", 
x"BCD141BDD000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BCD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BCD141BBD000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BCD111BCD000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"BCD141BDD000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DBCD1421DAAD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"DBCD1411DACD", 
x"D1D000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DBCD1441DADD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCD1121DBAD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"BC11BC000000", 
x"DBCD1141DBBD", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBCD1111DBCD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBCD1141DBDD", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"DBCD1411DCCD", 
x"CD11CD000000", 
x"DB11DB000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBC141DAC000", 
x"DBCD1421DDAD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"B1B000000000", 
x"DBC141DDC000", 
x"DBCD1411DDCD", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBC141DDC000", 
x"DBCD1441DDDD", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBDA2121ABAA", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDA2141ABBA", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"DBDA2141ABCA", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDA2111ABDA", 
x"DB11DB000000", 
x"DBD211ABD000", 
x"DBD211ABD000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BADA", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA121BAA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DA1411BCDA", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"BDA111BDA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"BDA121BAA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA141BBA000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDA141BCA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDA111BDA000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"DA11DA000000", 
x"DB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DA11DA000000", 
x"B1B000000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DBDA1411DADA", 
x"DB11DB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DBDA1121DBAA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDA1141DBBA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDA1141DBCA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDA1111DBDA", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBDA1421DCAA", 
x"DB21AB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBDA1411DCDA", 
x"DB11DB000000", 
x"DBD141DCD000", 
x"DBD141DCD000", 
x"DA11DA000000", 
x"DB21AB000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBDA1441DDCA", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DBDA1411DDDA", 
x"DB11DB000000", 
x"DBD141DDD000", 
x"DBD141DDD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDB2141AB3B", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDB2121ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDB2141AB3B", 
x"DBDB2141ABBB", 
x"DBDB2141AB3B", 
x"BD11BD000000", 
x"DB21AB000000", 
x"DBDB2141ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DBDB2111ABDB", 
x"DBD211ABD000", 
x"DBD211ABD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBDB1141DB3B", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"B1B000000000", 
x"B3DB1421BAAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"BD3B1241BACB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BADB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB121BAB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BDB141BCB000", 
x"BDB141B3B000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B3DB1421BCAB", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B3DB1441BCCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3DB1411BCDB", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD3B1141BDAB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD3B1141BDCB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B3DB1411BDDB", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDB2141AB3B", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB121BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"BDB141BBB000", 
x"BDB141B3B000", 
x"BD11BD000000", 
x"B1B000000000", 
x"BDB141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDB111BDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBDB1141DB3B", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DBD141DDD000", 
x"D1D000000000", 
x"DBDB1421DAAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDB2141AB3B", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"D1D000000000", 
x"DBDB1441DACB", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DBDB1411DADB", 
x"DBD141DAD000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBDB1121DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDB1141DB3B", 
x"DBDB1141DBBB", 
x"DBDB1141DB3B", 
x"DBDB1141DB3B", 
x"DB11DB000000", 
x"DBDB1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBDB1111DBDB", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"DBDB1421DCAB", 
x"D1D000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BDB141B3B000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DBDB1411DCDB", 
x"DBD141DCD000", 
x"DBD141DCD000", 
x"D1D000000000", 
x"DBDB1421DDAB", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBDB1141DB3B", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"DBDB1441DDCB", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DBD141DDD000", 
x"DBDB1411DDDB", 
x"DBD141DDD000", 
x"DBD141DDD000", 
x"000000000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDC2121ABAC", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDC2141ABBC", 
x"BD11BD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDC2141ABCC", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DB11DB000000", 
x"DBDC2111ABDC", 
x"DBD211ABD000", 
x"DC21AC000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DBD141DDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B3DC1411BADC", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B3DC1411BCDC", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC121BAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BBC000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDC141BCC000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BDC111BDC000", 
x"BD11BD000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DBD141DDD000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDC1421DAAC", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DBDC1441DACC", 
x"DC21AC000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBDC1411DADC", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDC1121DBAC", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDC1141DBBC", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDC1141DBCC", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBDC1111DBDC", 
x"DBD111DBD000", 
x"DC11DC000000", 
x"DB21AB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DB11DB000000", 
x"DBDC1411DCDC", 
x"DC11DC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBDC1421DDAC", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DBD141DDD000", 
x"DB11DB000000", 
x"DBDC1411DDDC", 
x"DBD141DDD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDD2121ABAD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBDD2141ABCD", 
x"DBD211ABD000", 
x"DB11DB000000", 
x"DBD211ABD000", 
x"DBDD2111ABDD", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"DB11DB000000", 
x"BDD121BAD000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"DB11DB000000", 
x"BDD141BCD000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"BDD111BDD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD121BAD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BDD141BCD000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BDD111BDD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBDD1421DAAD", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DBDD1441DACD", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DBD141DAD000", 
x"DBDD1411DADD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDD1121DBAD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDD1141DBBD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBDD1141DBCD", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBDD1111DBDD", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DBDD1421DCAD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DB11DB000000", 
x"DBD141DCD000", 
x"DBDD1411DCDD", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DD11DD000000", 
x"DBDD1411DDDD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DCA211ACA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DC11DC000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCAA2111ACAA", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCAA2141ACBA", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CA11CA000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAA2121ACDA", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DC11DC000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CAA111CAA000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"CAA121CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCAA1211DAAA", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCAA1241DABA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAA1221DADA", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCAA1411DBAA", 
x"DCA141DBA000", 
x"DC21AC000000", 
x"DCA141DBA000", 
x"DCAA1441DBBA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCAA1421DBDA", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCAA1111DCAA", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCAA1141DCBA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAA1121DCCA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAA1121DCDA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAA1411DDAA", 
x"DCA141DDA000", 
x"DC21AC000000", 
x"DCA141DDA000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"DCAB2211AAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"CAB211AAB000", 
x"DCA211ACA000", 
x"DCAB2221AACB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCAB2221AADB", 
x"DC11DC000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"DCA211ACA000", 
x"DCAB2111ACAB", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"CAB221ACB000", 
x"DCAB2141ACBB", 
x"CAB221ACB000", 
x"CAB221ACB000", 
x"CA11CA000000", 
x"DCAB2121ACCB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAB2121ACDB", 
x"DC11DC000000", 
x"DC21AC000000", 
x"DCA121DAA000", 
x"AB11AB000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"CAB221ADB000", 
x"DCA111DCA000", 
x"DCAB1141DC3B", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"CAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"DCA211ACA000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"B1B000000000", 
x"CAB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CAB121CDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCA111DCA000", 
x"DCAB1141DC3B", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"CA11CA000000", 
x"CAB211AAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA3B1141CACB", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA3B1141CADB", 
x"DC11DC000000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CAB141CBB000", 
x"CA11CA000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"DC11DC000000", 
x"AB21CB000000", 
x"CA11CA000000", 
x"CAB111CAB000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CAB121CCB000", 
x"CA11CA000000", 
x"CAB121CCB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"AB11AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"CAB121CDB000", 
x"DCA111DCA000", 
x"DCAB1141DC3B", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"AB21DB000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"DCAB1211DAAB", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"DCA211ACA000", 
x"DCAB1221DACB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCAB1221DADB", 
x"DC11DC000000", 
x"D1D000000000", 
x"AB21DB000000", 
x"DCAB1411DBAB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DCAB1441DBBB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"CA11CA000000", 
x"DCAB1421DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DCAB1421DBDB", 
x"DC11DC000000", 
x"AB21DB000000", 
x"DCA111DCA000", 
x"DCAB1111DCAB", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCAB1141DC3B", 
x"DCAB1141DCBB", 
x"DCAB1141DC3B", 
x"DCAB1141DC3B", 
x"DC11DC000000", 
x"DCAB1121DCCB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAB1121DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA121DAA000", 
x"DCAB1411DDAB", 
x"DC21AC000000", 
x"DCA141DDA000", 
x"AB21DB000000", 
x"DCAB1441DDBB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DCA111DCA000", 
x"DCAB1141DC3B", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"DCAB1421DDDB", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DCAC2211AAAC", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"CAC211AAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCAC2111ACAC", 
x"DCA211ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DCAC2141ACBC", 
x"AC11AC000000", 
x"CA11CA000000", 
x"AC11AC000000", 
x"DCAC2121ACCC", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DCAC2121ACDC", 
x"AC11AC000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"CAC211AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DC11DC000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAC111CAC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC141CBC000", 
x"C1C000000000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"CAC121CCC000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCA111DCA000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"CAC121CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCAC1211DAAC", 
x"DCA121DAA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCAC1241DABC", 
x"D1D000000000", 
x"DCA211ACA000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"DCA141DBA000", 
x"DCAC1411DBAC", 
x"DCA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCAC1441DBBC", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"DCAC1421DBCC", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCAC1111DCAC", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAC1141DCBC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAC1121DCCC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAC1121DCDC", 
x"DC11DC000000", 
x"DCA121DAA000", 
x"DCA141DDA000", 
x"DCAC1411DDAC", 
x"DCA141DDA000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"DCAC1441DDBC", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"DCAD2211AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CAD211AAD000", 
x"CAD211AAD000", 
x"DC11DC000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCAD2111ACAD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAD2141ACBD", 
x"CA11CA000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAD2121ACCD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DCAD2121ACDD", 
x"DCA121DAA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DC11DC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"CAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DC11DC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"CAD121CDD000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"DC21AC000000", 
x"AD11AD000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CAD141CBD000", 
x"DC11DC000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CAD111CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD141CBD000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"CAD121CCD000", 
x"DC11DC000000", 
x"CAD121CCD000", 
x"DCA121DAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"AD11AD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CAD121CDD000", 
x"CAD121CDD000", 
x"DC11DC000000", 
x"CAD121CDD000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCAD1211DAAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCAD1241DABD", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCAD1221DACD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DC11DC000000", 
x"AD11AD000000", 
x"DCA141DBA000", 
x"DCA141DBA000", 
x"DC21AC000000", 
x"DCAD1411DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCAD1441DBBD", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCAD1421DBDD", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCAD1111DCAD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAD1141DCBD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAD1121DCCD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCAD1121DCDD", 
x"DCA121DAA000", 
x"DCA141DDA000", 
x"DC21AC000000", 
x"DCAD1411DDAD", 
x"DCA141DBA000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCAD1441DDBD", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCA141DDA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCAD1421DDDD", 
x"A1A000000000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCBA2211AABA", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"CBA211ABA000", 
x"BA11BA000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DCBA2141ACAA", 
x"CB21AB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCBA2111ACBA", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCBA2141ACCA", 
x"CB11CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCBA2141ACDA", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DCB211ACB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"CBA141CAA000", 
x"DCB221AAB000", 
x"CBA141CAA000", 
x"CBA141CAA000", 
x"CBA211ABA000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CAA000", 
x"CB21AB000000", 
x"CBA141CCA000", 
x"CBA141CCA000", 
x"CBA111CBA000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBA141CCA000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CBA141CDA000", 
x"DCB121DAB000", 
x"CBA141CDA000", 
x"CBA141CDA000", 
x"BA11BA000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCBA1241DAAA", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCBA1211DABA", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCBA1241DADA", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DCBA1411DBBA", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCBA1141DCAA", 
x"DC3B1141DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCBA1111DCBA", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCBA1141DCCA", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCBA1141DCDA", 
x"DC3B1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCBA1441DDAA", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCBA1411DDBA", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCBA1441DDDA", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DCBB2211AABB", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB3B2141ABAB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CBB211ABB000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB3B2141ABDB", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"DCBB2141ACAB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DCBB2111ACBB", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"CB11CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCBB2141ACDB", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"CBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CBB141CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBB141CDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"BB11BB000000", 
x"B3B141BDB000", 
x"B3B141BDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"CBB211ABB000", 
x"CBB141CAB000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB3B1141CBAB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB3B1141CBCB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB3B1141CBDB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBB141CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CBB111CBB000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBB141CDB000", 
x"BB11BB000000", 
x"CBB141CDB000", 
x"CBB141CDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCBB1241DAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCBB1211DABB", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCBB1241DADB", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"DCBB1411DBBB", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCBB1141DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCBB1111DCBB", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DCBB1141DCCB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCBB1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DCBB1411DDBB", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCBC2211AABC", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BC11BC000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB11CB000000", 
x"CBC211ABC000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"CB21AB000000", 
x"DCBC2141ACAC", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCBC2111ACBC", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"CB11CB000000", 
x"DCBC2141ACCC", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DCBC2141ACDC", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBC211ABC000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"DCB211ACB000", 
x"CBC141CAC000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CBC141CAC000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBC111CBC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CB11CB000000", 
x"CBC141CCC000", 
x"CBC141CCC000", 
x"C1C000000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"BC11BC000000", 
x"B1B000000000", 
x"CBC141CDC000", 
x"DCB111DCB000", 
x"CBC141CDC000", 
x"CBC141CDC000", 
x"C1C000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DCBC1241DAAC", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCBC1211DABC", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DCBC1241DACC", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCBC1411DBBC", 
x"DCB141DBB000", 
x"BC11BC000000", 
x"CB11CB000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"DCBC1141DCAC", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCBC1111DCBC", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DCBC1141DCCC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC3B1141DCDB", 
x"DCBC1141DCDC", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCBC1441DDAC", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCBC1411DDBC", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCBD2211AABD", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"BD11BD000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"CBD211ABD000", 
x"DC21AC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"DCBD2141ACAD", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCBD2111ACBD", 
x"DC21AC000000", 
x"CB11CB000000", 
x"DC21AC000000", 
x"DCBD2141ACCD", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCBD2141ACDD", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CBD211ABD000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DCB121DAB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DCB111DCB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"C1C000000000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CBD211ABD000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"CBD141CAD000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CBD111CBD000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CBD141CCD000", 
x"CBD141CCD000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CBD141CDD000", 
x"C1C000000000", 
x"DCB121DAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CBD141CDD000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"CBD141CDD000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DC21AC000000", 
x"DCBD1241DAAD", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCBD1211DABD", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCBD1241DADD", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCBD1411DBBD", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"DC11DC000000", 
x"DCBD1141DCAD", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCBD1111DCBD", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DC11DC000000", 
x"DCBD1141DCCD", 
x"DC11DC000000", 
x"DC3B1141DCDB", 
x"DC11DC000000", 
x"DCBD1141DCDD", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DC21AC000000", 
x"DCBD1441DDAD", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DCBD1411DDBD", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCB141DDB000", 
x"DC11DC000000", 
x"DCBD1441DDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCCA2211AACA", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"CCA211ACA000", 
x"DCCA2141ACBA", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCA2111ACCA", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCCA2141ACDA", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CCA211ACA000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DCC211ACC000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DC11DC000000", 
x"CA11CA000000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"CCA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA111CCA000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCA141CDA000", 
x"CCA141CDA000", 
x"DCC121DAC000", 
x"CCA141CDA000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC141DBC000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"DCCA1221DAAA", 
x"D1D000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCCA1241DABA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCCA1211DACA", 
x"DCC121DAC000", 
x"DCC211ACC000", 
x"DCC121DAC000", 
x"DCCA1241DADA", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCCA1421DBAA", 
x"D1D000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCCA1411DBCA", 
x"DCC141DBC000", 
x"CC11CC000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCCA1121DCAA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCA1141DCBA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCA1111DCCA", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCCA1141DCDA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCA1421DDAA", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DCCA1411DDCA", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DCCA1441DDDA", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"DCCB2221AAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"CCB221AAB000", 
x"DC21AC000000", 
x"DCCB2211AACB", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"DCCB2121ACAB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"CCB211ACB000", 
x"DCC211ACC000", 
x"DCCB2111ACCB", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"DCCB2141ACDB", 
x"DC11DC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB211ACB000", 
x"DCC211ACC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CCB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"B1B000000000", 
x"CCB141CDB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCC121DAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CCB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"CCB121CAB000", 
x"C1C000000000", 
x"CCB211ACB000", 
x"DCC211ACC000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CC11CC000000", 
x"CCB121CAB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CCB111CCB000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC3B1141CCDB", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"DCC121DAC000", 
x"C1C000000000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"CCB141CDB000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCCB1221DAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"CB21AB000000", 
x"DCCB1241DABB", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DCC121DAC000", 
x"DCCB1211DACB", 
x"DCC211ACC000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"DCCB1241DADB", 
x"DC11DC000000", 
x"D1D000000000", 
x"B1B000000000", 
x"DCCB1421DBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCCB1411DBCB", 
x"CC11CC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCCB1121DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"CB11CB000000", 
x"DCCB1141DCBB", 
x"CB11CB000000", 
x"CB11CB000000", 
x"DCC111DCC000", 
x"DCCB1111DCCB", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DCCB1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCCB1421DDAB", 
x"DCC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCCB1411DDCB", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCCB1441DDDB", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCC2121ACAC", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCC2141ACBC", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCCC2111ACCC", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCC2141ACDC", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC121CAC000", 
x"CCC121CAC000", 
x"DCC211ACC000", 
x"CCC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCC141CBC000", 
x"CCC141CBC000", 
x"CC11CC000000", 
x"CCC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CCC111CCC000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC121DAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC141DBC000", 
x"C1C000000000", 
x"CCC141CDC000", 
x"CCC141CDC000", 
x"DCC111DCC000", 
x"CCC141CDC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCCC1221DAAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCCC1241DABC", 
x"D1D000000000", 
x"DCC121DAC000", 
x"DCC121DAC000", 
x"DCCC1211DACC", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCCC1421DBAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"DCC141DBC000", 
x"DCCC1411DBCC", 
x"DCC141DBC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCC1121DCAC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCC1141DCBC", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCCC1111DCCC", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCC1141DCDC", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DCCD2211AACD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCD2121ACAD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCCD2141ACBD", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCCD2111ACCD", 
x"CCD211ACD000", 
x"CCD211ACD000", 
x"DC11DC000000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"CCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC211ACC000", 
x"CCD211ACD000", 
x"CCD121CAD000", 
x"CCD121CAD000", 
x"DC11DC000000", 
x"CCD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CD11CD000000", 
x"CCD141CBD000", 
x"CCD141CBD000", 
x"DC11DC000000", 
x"CCD141CBD000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CCD111CCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DCC121DAC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCCD1221DAAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCCD1241DABD", 
x"DCC121DAC000", 
x"DCC121DAC000", 
x"DCC211ACC000", 
x"DCCD1211DACD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCCD1241DADD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCCD1421DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"DCC141DBC000", 
x"CC11CC000000", 
x"DCCD1411DBCD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCD1121DCAD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCD1141DCBD", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCCD1111DCCD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCCD1141DCDD", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC121DAC000", 
x"DCCD1421DDAD", 
x"D1D000000000", 
x"D1D000000000", 
x"DCC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DCCD1411DDCD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCCD1441DDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"DCDA2211AADA", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DCDA2121ACAA", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDA2141ACBA", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDA2141ACCA", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CD11CD000000", 
x"DCDA2111ACDA", 
x"DCD211ACD000", 
x"DC11DC000000", 
x"DCD211ACD000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"CDA211ADA000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"CDA211ADA000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"CDA121CAA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCD211ACD000", 
x"CDA211ADA000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"CDA121CAA000", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"CDA141CCA000", 
x"CDA141CBA000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDA141CCA000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CDA111CDA000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DCD211ACD000", 
x"DCDA1211DADA", 
x"DCD121DAD000", 
x"DC11DC000000", 
x"DCD121DAD000", 
x"DCDA1421DBAA", 
x"D1D000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"DCDA1441DBBA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCDA1411DBDA", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DCD141DBD000", 
x"DCDA1121DCAA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDA1141DCBA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDA1141DCCA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDA1111DCDA", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DCD121DAD000", 
x"DCDA1441DDBA", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCDA1411DDDA", 
x"DCD141DDD000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"000000000000", 
x"DCDB2221AAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"CDB221AAB000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"DCDB2211AADB", 
x"DC11DC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"CD11CD000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"DCDB2121ACAB", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DCDB2141ACBB", 
x"B1B000000000", 
x"B1B000000000", 
x"DC21AC000000", 
x"DCDB2141ACCB", 
x"DC21AC000000", 
x"CD11CD000000", 
x"DCD211ACD000", 
x"DCDB2111ACDB", 
x"DC11DC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"CDB211ADB000", 
x"DC11DC000000", 
x"DCDB1141DC3B", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCD211ACD000", 
x"B1B000000000", 
x"CDB211ADB000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB121CAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CCB000", 
x"B1B000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DCDB1141DC3B", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DCD211ACD000", 
x"C1C000000000", 
x"CDB211ADB000", 
x"DC11DC000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"CDB141CBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CD11CD000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"CDB121CAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"CDB141CBB000", 
x"CDB141CCB000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CDB141CCB000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD3B1141CDAB", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"CDB111CDB000", 
x"DC11DC000000", 
x"DCDB1141DC3B", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CD11CD000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"DCDB1221DAAB", 
x"DC21AC000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DCDB1241DABB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DC21AC000000", 
x"DCDB1241DACB", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"DCD121DAD000", 
x"DCDB1211DADB", 
x"DC11DC000000", 
x"DCD121DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DCDB1411DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DCDB1121DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDB1141DC3B", 
x"DCDB1141DCBB", 
x"DCDB1141DC3B", 
x"DCDB1141DC3B", 
x"DC11DC000000", 
x"DCDB1141DCCB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCDB1111DCDB", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"DCDB1421DDAB", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DC11DC000000", 
x"DCDB1141DC3B", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD141DDD000", 
x"DCDB1411DDDB", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDC2121ACAC", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDC2141ACBC", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDC2141ACCC", 
x"CD11CD000000", 
x"DCD211ACD000", 
x"DCD211ACD000", 
x"DCDC2111ACDC", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCD141DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC121CAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDC141CBC000", 
x"C1C000000000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CDC141CCC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CDC111CDC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1221DAAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1241DABC", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDC1241DACC", 
x"DCD211ACD000", 
x"DCD121DAD000", 
x"DCD121DAD000", 
x"DCDC1211DADC", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1421DBAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1441DBBC", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCD141DBD000", 
x"DCD141DBD000", 
x"DCDC1411DBDC", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDC1121DCAC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDC1141DCBC", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDC1141DCCC", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCDC1111DCDC", 
x"DCD111DCD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1421DDAC", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DCDC1441DDBC", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DCD141DDD000", 
x"DCD141DDD000", 
x"DCDC1411DDDC", 
x"DCD141DDD000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DCDD2211AADD", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDD2121ACAD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCDD2141ACBD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CD11CD000000", 
x"DCD211ACD000", 
x"DCD211ACD000", 
x"DC11DC000000", 
x"DCDD2111ACDD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CDD211ADD000", 
x"CDD211ADD000", 
x"DC11DC000000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"CDD211ADD000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCD211ACD000", 
x"CDD121CAD000", 
x"CDD121CAD000", 
x"DC11DC000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CDD141CBD000", 
x"CDD141CBD000", 
x"DC11DC000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD121CAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CDD141CBD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CDD111CDD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"CDD111CDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCDD1221DAAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCDD1241DABD", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"DCD121DAD000", 
x"DCD121DAD000", 
x"DC11DC000000", 
x"DCDD1211DADD", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DCDD1421DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DCDD1441DBBD", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"DCD141DBD000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DCDD1411DBDD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDD1121DCAD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDD1141DCBD", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCDD1141DCCD", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCDD1111DCDD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DCD121DAD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DCDD1411DDDD", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DDA211ADA000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDAA2111ADAA", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAA2121ADCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AA11AA000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAA121DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DAA111DAA000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DD11DD000000", 
x"DDAA1411DBAA", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDAA1441DBBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAA1421DBCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDAA1411DCAA", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DAA121DCA000", 
x"DDAA1441DCBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAA1421DCCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDAA1111DDAA", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDAA1141DDBA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDAA1121DDCA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"DDAB2211AAAB", 
x"A1A000000000", 
x"D1D000000000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"DDAB2221AACB", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"DDAB2221AADB", 
x"D1D000000000", 
x"DD11DD000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA211ADA000", 
x"DDAB2111ADAB", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DAB221ADB000", 
x"DDAB2141ADBB", 
x"DAB221ADB000", 
x"DAB221ADB000", 
x"DDA141DCA000", 
x"DDAB2121ADCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DDAB2121ADDB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DAB211AAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"AB11AB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB111DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DAB121DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDA111DDA000", 
x"DAB121DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DAB211AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"DAB221ACB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"DAB221ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"AB21CB000000", 
x"AB11AB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB11AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"AB21CB000000", 
x"A1A000000000", 
x"AB21CB000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DDA141DCA000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDA111DDA000", 
x"DAB121DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DDAB1211DAAB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DAB111DAB000", 
x"DA11DA000000", 
x"DDAB1221DACB", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDAB1221DADB", 
x"DA11DA000000", 
x"DD11DD000000", 
x"AB21DB000000", 
x"DDAB1411DBAB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"DAB141DBB000", 
x"AB21DB000000", 
x"DDAB1421DBCB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DDAB1421DBDB", 
x"AB21DB000000", 
x"AB21DB000000", 
x"DDA141DCA000", 
x"DDAB1411DCAB", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"DAB121DCB000", 
x"D1D000000000", 
x"DDAB1421DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"DDAB1421DCDB", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDAB1111DDAB", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DAB121DDB000", 
x"DDAB1141DDBB", 
x"DAB121DDB000", 
x"DAB121DDB000", 
x"DD11DD000000", 
x"DDAB1121DDCB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDAB1121DDDB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DDAC2211AAAC", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DAC211AAC000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"DDAC2221AADC", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"DD11DD000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDAC2111ADAC", 
x"DDA211ADA000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"DDAC2141ADBC", 
x"D1D000000000", 
x"DDA141DCA000", 
x"DAC221ADC000", 
x"DDAC2121ADCC", 
x"DAC221ADC000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DDAC2121ADDC", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAC211AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"DAC221ADC000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AC11AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"AC21DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"DAC141DBC000", 
x"D1D000000000", 
x"DDA141DCA000", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"AC21DC000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DAC121DDC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DAC211AAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"AC11AC000000", 
x"DDA211ADA000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"AC11AC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DA11DA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DDA141DBA000", 
x"C1C000000000", 
x"DAC141DBC000", 
x"C1C000000000", 
x"DDA141DCA000", 
x"C1C000000000", 
x"DAC121DCC000", 
x"C1C000000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DAC121DDC000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDAC1211DAAC", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDAC1241DABC", 
x"DA11DA000000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DAC111DAC000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDAC1221DADC", 
x"DD11DD000000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDAC1411DBAC", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAC1441DBBC", 
x"D1D000000000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DAC141DBC000", 
x"DA11DA000000", 
x"D1D000000000", 
x"DDAC1421DBDC", 
x"DD11DD000000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDAC1411DCAC", 
x"DDA141DCA000", 
x"AC21DC000000", 
x"AC21DC000000", 
x"DDAC1441DCBC", 
x"AC21DC000000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DAC121DCC000", 
x"DA11DA000000", 
x"AC21DC000000", 
x"DDAC1421DCDC", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDAC1111DDAC", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDAC1141DDBC", 
x"DD11DD000000", 
x"DAC121DDC000", 
x"DAC121DDC000", 
x"DDAC1121DDCC", 
x"DAC121DDC000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DDAC1121DDDC", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DDAD2211AAAD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"DAD211AAD000", 
x"DAD211AAD000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDAD2111ADAD", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"DDA141DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DAD211AAD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"AD11AD000000", 
x"AD11AD000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"AD11AD000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD141DBD000", 
x"DDA141DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DAD121DCD000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDAD1211DAAD", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DAD111DAD000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDAD1411DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAD1441DBBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAD1421DBCD", 
x"DA11DA000000", 
x"DAD141DBD000", 
x"DAD141DBD000", 
x"DD11DD000000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDAD1411DCAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAD1441DCBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDAD1421DCCD", 
x"DA11DA000000", 
x"DAD121DCD000", 
x"DAD121DCD000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDAD1111DDAD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDAD1141DDBD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDAD1121DDCD", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDAD1121DDDD", 
x"A1A000000000", 
x"DDB221AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDBA2211AABA", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"DBA211ABA000", 
x"BA11BA000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDBA2141ADAA", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDBA2111ADBA", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDBA2141ADCA", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"DDB211ADB000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DDB221AAB000", 
x"A1A000000000", 
x"D1D000000000", 
x"DBA211ABA000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"DB21AB000000", 
x"A1A000000000", 
x"D1D000000000", 
x"BA11BA000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"A1A000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DBA141DAA000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBA111DBA000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DBA141DAA000", 
x"DDB221AAB000", 
x"DBA141DAA000", 
x"DBA141DAA000", 
x"DDBA1211DABA", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDBA1241DACA", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDBA1241DADA", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DBA111DBA000", 
x"DDBA1411DBBA", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBA141DCA000", 
x"DB21AB000000", 
x"DBA141DCA000", 
x"DBA141DCA000", 
x"DDBA1411DCBA", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDBA1441DCDA", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDBA1141DDAA", 
x"DDB121DAB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDBA1111DDBA", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDBA1141DDCA", 
x"DDB141DCB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDBA1141DDDA", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"DDB221AAB000", 
x"000000000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"DDBB2211AABB", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DB3B2141ABAB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB3B2141ABCB", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"DDBB2111ADBB", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"DBB211ABB000", 
x"B3B141BAB000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"BB11BB000000", 
x"B3B141BCB000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"DDB221AAB000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DBB211ABB000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B3B141BAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B3B141BCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"BB11BB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDBB1241DAAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDBB1211DABB", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"DDBB1241DACB", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB3B1141DBAB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DBB111DBB000", 
x"DB11DB000000", 
x"DB3B1141DBCB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB3B1141DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DDBB1441DCAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"DDBB1411DCBB", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDBB1141DDAB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDBB1111DDBB", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDBB1141DDCB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"000000000000", 
x"DDB221AAB000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDBC2211AABC", 
x"DDB221AAB000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"C1C000000000", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BC11BC000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDBC2141ADAC", 
x"D1D000000000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDBC2111ADBC", 
x"DDB211ADB000", 
x"C1C000000000", 
x"DDB141DCB000", 
x"DDBC2141ADCC", 
x"C1C000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDBC2141ADDC", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBC211ABC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DDB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBC211ABC000", 
x"DB21AB000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDB211ADB000", 
x"C1C000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BC11BC000000", 
x"B1B000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"DDB121DAB000", 
x"DBC141DAC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DDB141DCB000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DBC141DDC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"DDBC1241DAAC", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDBC1211DABC", 
x"DDB121DAB000", 
x"DBC141DAC000", 
x"B1B000000000", 
x"DBC141DAC000", 
x"DBC141DAC000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"DDBC1241DADC", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DDBC1411DBBC", 
x"DB11DB000000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DBC111DBC000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"C1C000000000", 
x"DB21AB000000", 
x"DDBC1441DCAC", 
x"C1C000000000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDBC1411DCBC", 
x"DDB141DCB000", 
x"DBC141DCC000", 
x"B1B000000000", 
x"DBC141DCC000", 
x"DBC141DCC000", 
x"C1C000000000", 
x"DB11DB000000", 
x"DDBC1441DCDC", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB121DAB000", 
x"DDBC1141DDAC", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDBC1111DDBC", 
x"DDB111DDB000", 
x"DBC141DDC000", 
x"DDB141DCB000", 
x"DDBC1141DDCC", 
x"DBC141DDC000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDBC1141DDDC", 
x"DD11DD000000", 
x"000000000000", 
x"DDB221AAB000", 
x"000000000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDBD2211AABD", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"BD11BD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"DB11DB000000", 
x"DBD211ABD000", 
x"DBD211ABD000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"DDBD2141ADAD", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDBD2111ADBD", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"DDBD2141ADCD", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DBD211ABD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DDB121DAB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"DDB111DDB000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DDB221AAB000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DBD211ABD000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"DB11DB000000", 
x"BD11BD000000", 
x"BD11BD000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"BD11BD000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"DBD141DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"D1D000000000", 
x"DDBD1241DAAD", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDBD1211DABD", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"DDBD1241DACD", 
x"DBD141DAD000", 
x"DDB211ADB000", 
x"DBD141DAD000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DDBD1411DBBD", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"DBD111DBD000", 
x"D1D000000000", 
x"DB21AB000000", 
x"D1D000000000", 
x"DDBD1441DCAD", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDBD1411DCBD", 
x"D1D000000000", 
x"B1B000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DBD141DCD000", 
x"DB11DB000000", 
x"DBD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB121DAB000", 
x"DD11DD000000", 
x"DDBD1141DDAD", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDBD1111DDBD", 
x"DD11DD000000", 
x"DDB141DCB000", 
x"DD11DD000000", 
x"DDBD1141DDCD", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDBD1141DDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDCA2211AACA", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CA11CA000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DDCA2121ADAA", 
x"D1D000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"DDCA2141ADBA", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DDCA2111ADCA", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DCA211ACA000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DCA121DAA000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"DCA141DBA000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"DDC211ADC000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CA11CA000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DCA121DAA000", 
x"C1C000000000", 
x"DDC121DAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC141DBC000", 
x"C1C000000000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DCA121DAA000", 
x"DDCA1241DABA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDCA1211DACA", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDCA1241DADA", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"DDCA1421DBAA", 
x"DCA141DBA000", 
x"DC21AC000000", 
x"DCA141DBA000", 
x"DDCA1441DBBA", 
x"D1D000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDCA1411DBCA", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDCA1441DBDA", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DCA111DCA000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DDCA1411DCCA", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DDCA1121DDAA", 
x"DD11DD000000", 
x"DDC121DAC000", 
x"DD11DD000000", 
x"DDCA1141DDBA", 
x"DD11DD000000", 
x"DDC141DBC000", 
x"DD11DD000000", 
x"DDCA1111DDCA", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDCA1141DDDA", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"DDCB2221AAAB", 
x"DDC221AAC000", 
x"D1D000000000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DCB221AAB000", 
x"DDC221AAC000", 
x"DDCB2211AACB", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB11CB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"DC11DC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"CB21AB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DCB211ACB000", 
x"DC21AC000000", 
x"CB11CB000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDCB2121ADAB", 
x"DDC121DAC000", 
x"D1D000000000", 
x"B1B000000000", 
x"DDCB2141ADBB", 
x"B1B000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DDCB2111ADCB", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"DDCB2141ADDB", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB211ACB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"CB11CB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB121DAB000", 
x"DDC121DAC000", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"B1B000000000", 
x"DCB141DDB000", 
x"DDC111DDC000", 
x"B1B000000000", 
x"C1C000000000", 
x"DCB221AAB000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"DCB211ACB000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB21AB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"CB11CB000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"DCB121DAB000", 
x"DDC121DAC000", 
x"C1C000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DCB141DDB000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDCB1221DAAB", 
x"DDC221AAC000", 
x"D1D000000000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DCB121DAB000", 
x"DDC121DAC000", 
x"DDCB1211DACB", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"DDCB1241DADB", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"B1B000000000", 
x"DDCB1421DBAB", 
x"B1B000000000", 
x"B1B000000000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"DCB141DBB000", 
x"B1B000000000", 
x"DDCB1411DBCB", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDCB1441DBDB", 
x"DC11DC000000", 
x"B1B000000000", 
x"DC11DC000000", 
x"DC3B1141DCAB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DCB111DCB000", 
x"DC11DC000000", 
x"DDCB1411DCCB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC3B1141DCDB", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DDCB1121DDAB", 
x"DDC121DAC000", 
x"DD11DD000000", 
x"DCB141DDB000", 
x"DDCB1141DDBB", 
x"DCB141DDB000", 
x"DCB141DDB000", 
x"DDC111DDC000", 
x"DDCB1111DDCB", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"DDCB1141DDDB", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDCC2211AACC", 
x"DDC221AAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDCC2111ADCC", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCC211ACC000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCC211ACC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"CC11CC000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC121DAC000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC141DBC000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDCC1221DAAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDCC1241DABC", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDCC1211DACC", 
x"DDC121DAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDCC1421DBAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDCC1441DBBC", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDCC1411DBCC", 
x"DDC141DBC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DCC111DCC000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDCC1121DDAC", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDCC1141DDBC", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDCC1111DDCC", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDCD2211AACD", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"CD11CD000000", 
x"DCD211ACD000", 
x"DCD211ACD000", 
x"DC11DC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DDCD2121ADAD", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDCD2141ADBD", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDCD2111ADCD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DCD211ACD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DCD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DCD211ACD000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DDC121DAC000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DCD111DCD000", 
x"CD11CD000000", 
x"CD11CD000000", 
x"DDC111DDC000", 
x"CD11CD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC221AAC000", 
x"DDCD1221DAAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DDCD1241DABD", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDCD1211DACD", 
x"DCD121DAD000", 
x"DCD121DAD000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DDCD1421DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"DDCD1441DBBD", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDCD1411DBCD", 
x"DCD141DBD000", 
x"DCD141DBD000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DDCD1411DCCD", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DCD111DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC121DAC000", 
x"DDCD1121DDAD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC141DBC000", 
x"DDCD1141DDBD", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDCD1111DDCD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDCD1141DDDD", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDDA2211AADA", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDA211ADA000", 
x"DDD121DAD000", 
x"DDDA2141ADBA", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"DDDA2141ADCA", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DDDA2111ADDA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDD121DAD000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"DDA141DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"DDA211ADA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"A1A000000000", 
x"A1A000000000", 
x"A1A000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"A1A000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"DA11DA000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDD121DAD000", 
x"DDA141DBA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"DDA141DCA000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DDA111DDA000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DA11DA000000", 
x"DDDA1211DADA", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"DD11DD000000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDA141DBA000", 
x"DDDA1441DBBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDA1441DBCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDA1411DBDA", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DD11DD000000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDA141DCA000", 
x"DDDA1441DCBA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDA1441DCCA", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDA1411DCDA", 
x"DDD141DCD000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDA111DDA000", 
x"DDDA1141DDBA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDA1141DDCA", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDA1111DDDA", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"000000000000", 
x"DDDB2221AAAB", 
x"000000000000", 
x"D1D000000000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"DDB221AAB000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDB2211AADB", 
x"D1D000000000", 
x"DD11DD000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB11DB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDDB2121ADAB", 
x"D1D000000000", 
x"DDD121DAD000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DDDB2141ADCB", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DDDB2111ADDB", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB211ADB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB121DAB000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"DDB141DCB000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DDB111DDB000", 
x"B1B000000000", 
x"DDD111DDD000", 
x"000000000000", 
x"DDB221AAB000", 
x"000000000000", 
x"D1D000000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"DB21AB000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB211ADB000", 
x"D1D000000000", 
x"DD11DD000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"DB11DB000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"DB21AB000000", 
x"000000000000", 
x"D1D000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"B1B000000000", 
x"000000000000", 
x"B1B000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"D1D000000000", 
x"DDDB1221DAAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"DDB121DAB000", 
x"D1D000000000", 
x"DDDB1241DACB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"DDDB1211DADB", 
x"DDD121DAD000", 
x"DD11DD000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DB11DB000000", 
x"DDDB1411DBDB", 
x"DB11DB000000", 
x"DB11DB000000", 
x"D1D000000000", 
x"DDDB1421DCAB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"DDB141DCB000", 
x"D1D000000000", 
x"DDDB1441DCCB", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DDDB1411DCDB", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDB1121DDAB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DDB111DDB000", 
x"DD11DD000000", 
x"DDDB1141DDCB", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"DDDB1111DDDB", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"000000000000", 
x"000000000000", 
x"DDDC2221AAAC", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC2211AADC", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC2121ADAC", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC2141ADBC", 
x"DDD141DBD000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDC2111ADDC", 
x"DDD111DDD000", 
x"000000000000", 
x"000000000000", 
x"DDC221AAC000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"DC21AC000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDD111DDD000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC211ADC000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC121DAC000", 
x"DDD121DAD000", 
x"C1C000000000", 
x"C1C000000000", 
x"DDC141DBC000", 
x"DDD141DBD000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDD111DDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC1221DAAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC1241DABC", 
x"D1D000000000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDC121DAC000", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"DDDC1211DADC", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC1421DBAC", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDC1441DBBC", 
x"D1D000000000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDC141DBC000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DDDC1411DBDC", 
x"DD11DD000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DC11DC000000", 
x"DDDC1411DCDC", 
x"DC11DC000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDC1121DDAC", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDC1141DDBC", 
x"DD11DD000000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDC111DDC000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDDC1111DDDC", 
x"DDD111DDD000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"000000000000", 
x"000000000000", 
x"000000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DD11DD000000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD121DAD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DBD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDD141DCD000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDD111DDD000", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1221DAAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1241DABD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1241DACD", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"DDD121DAD000", 
x"DDDD1211DADD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1421DBAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1441DBBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1441DBCD", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DDD141DBD000", 
x"DDDD1411DBDD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1421DCAD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1441DCBD", 
x"D1D000000000", 
x"D1D000000000", 
x"D1D000000000", 
x"DDDD1441DCCD", 
x"DDD141DCD000", 
x"DDD141DCD000", 
x"DDD141DCD000", 
x"DDDD1411DCDD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDD1121DDAD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDD1141DDBD", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DD11DD000000", 
x"DDDD1141DDCD", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDD111DDD000", 
x"DDDD1111DDDD");
begin
process(clk)
begin
if (clk'event and clk='1') then
data <= memory(to_integer(unsigned(addr)));
end if;
end process;
end Behavioral;

